magic
tech sky130A
magscale 1 2
timestamp 1651151325
<< obsli1 >>
rect 1104 2159 54096 54961
<< obsm1 >>
rect 14 2128 54910 54992
<< metal2 >>
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16302 0 16358 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27250 0 27306 800
rect 27802 0 27858 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29274 0 29330 800
rect 29826 0 29882 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 33966 0 34022 800
rect 34518 0 34574 800
rect 35070 0 35126 800
rect 35530 0 35586 800
rect 36082 0 36138 800
rect 36634 0 36690 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43350 0 43406 800
rect 43902 0 43958 800
rect 44454 0 44510 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54850 0 54906 800
<< obsm2 >>
rect 20 856 54904 54992
rect 20 734 146 856
rect 314 734 606 856
rect 774 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2170 856
rect 2338 734 2722 856
rect 2890 734 3182 856
rect 3350 734 3734 856
rect 3902 734 4286 856
rect 4454 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5850 856
rect 6018 734 6310 856
rect 6478 734 6862 856
rect 7030 734 7414 856
rect 7582 734 7874 856
rect 8042 734 8426 856
rect 8594 734 8978 856
rect 9146 734 9438 856
rect 9606 734 9990 856
rect 10158 734 10542 856
rect 10710 734 11002 856
rect 11170 734 11554 856
rect 11722 734 12106 856
rect 12274 734 12566 856
rect 12734 734 13118 856
rect 13286 734 13670 856
rect 13838 734 14130 856
rect 14298 734 14682 856
rect 14850 734 15234 856
rect 15402 734 15694 856
rect 15862 734 16246 856
rect 16414 734 16798 856
rect 16966 734 17258 856
rect 17426 734 17810 856
rect 17978 734 18362 856
rect 18530 734 18822 856
rect 18990 734 19374 856
rect 19542 734 19926 856
rect 20094 734 20386 856
rect 20554 734 20938 856
rect 21106 734 21490 856
rect 21658 734 21950 856
rect 22118 734 22502 856
rect 22670 734 23054 856
rect 23222 734 23514 856
rect 23682 734 24066 856
rect 24234 734 24618 856
rect 24786 734 25078 856
rect 25246 734 25630 856
rect 25798 734 26182 856
rect 26350 734 26642 856
rect 26810 734 27194 856
rect 27362 734 27746 856
rect 27914 734 28206 856
rect 28374 734 28758 856
rect 28926 734 29218 856
rect 29386 734 29770 856
rect 29938 734 30322 856
rect 30490 734 30782 856
rect 30950 734 31334 856
rect 31502 734 31886 856
rect 32054 734 32346 856
rect 32514 734 32898 856
rect 33066 734 33450 856
rect 33618 734 33910 856
rect 34078 734 34462 856
rect 34630 734 35014 856
rect 35182 734 35474 856
rect 35642 734 36026 856
rect 36194 734 36578 856
rect 36746 734 37038 856
rect 37206 734 37590 856
rect 37758 734 38142 856
rect 38310 734 38602 856
rect 38770 734 39154 856
rect 39322 734 39706 856
rect 39874 734 40166 856
rect 40334 734 40718 856
rect 40886 734 41270 856
rect 41438 734 41730 856
rect 41898 734 42282 856
rect 42450 734 42834 856
rect 43002 734 43294 856
rect 43462 734 43846 856
rect 44014 734 44398 856
rect 44566 734 44858 856
rect 45026 734 45410 856
rect 45578 734 45962 856
rect 46130 734 46422 856
rect 46590 734 46974 856
rect 47142 734 47526 856
rect 47694 734 47986 856
rect 48154 734 48538 856
rect 48706 734 49090 856
rect 49258 734 49550 856
rect 49718 734 50102 856
rect 50270 734 50654 856
rect 50822 734 51114 856
rect 51282 734 51666 856
rect 51834 734 52218 856
rect 52386 734 52678 856
rect 52846 734 53230 856
rect 53398 734 53782 856
rect 53950 734 54242 856
rect 54410 734 54794 856
<< obsm3 >>
rect 4208 2143 50608 54977
<< metal4 >>
rect 4208 2128 4528 54992
rect 19568 2128 19888 54992
rect 34928 2128 35248 54992
rect 50288 2128 50608 54992
<< labels >>
rlabel metal4 s 19568 2128 19888 54992 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 54992 6 VGND
port 1 nsew ground input
rlabel metal4 s 4208 2128 4528 54992 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 54992 6 VPWR
port 2 nsew power input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 4 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 5 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[0]
port 6 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[10]
port 7 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[11]
port 8 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[12]
port 9 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[13]
port 10 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[14]
port 11 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[15]
port 12 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[16]
port 13 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[17]
port 14 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[18]
port 15 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_adr_i[19]
port 16 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[1]
port 17 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[20]
port 18 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[21]
port 19 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[22]
port 20 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[23]
port 21 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[24]
port 22 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[25]
port 23 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_adr_i[26]
port 24 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[27]
port 25 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_adr_i[28]
port 26 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_adr_i[29]
port 27 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[2]
port 28 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[30]
port 29 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_adr_i[31]
port 30 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[3]
port 31 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[4]
port 32 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[5]
port 33 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[6]
port 34 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[7]
port 35 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[8]
port 36 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[9]
port 37 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 38 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[0]
port 39 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[10]
port 40 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[11]
port 41 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[12]
port 42 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[13]
port 43 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[14]
port 44 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[15]
port 45 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[16]
port 46 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[17]
port 47 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[18]
port 48 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[19]
port 49 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[1]
port 50 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[20]
port 51 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[21]
port 52 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[22]
port 53 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[23]
port 54 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[24]
port 55 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[25]
port 56 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_i[26]
port 57 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[27]
port 58 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[28]
port 59 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[29]
port 60 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[2]
port 61 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[30]
port 62 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[31]
port 63 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[3]
port 64 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[4]
port 65 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[5]
port 66 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[6]
port 67 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[7]
port 68 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[8]
port 69 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[9]
port 70 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[0]
port 71 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[10]
port 72 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[11]
port 73 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[12]
port 74 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[13]
port 75 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[14]
port 76 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_o[15]
port 77 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[16]
port 78 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[17]
port 79 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[18]
port 80 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[19]
port 81 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[1]
port 82 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_o[20]
port 83 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[21]
port 84 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_o[22]
port 85 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_o[23]
port 86 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[24]
port 87 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[25]
port 88 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_o[26]
port 89 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[27]
port 90 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_o[28]
port 91 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[29]
port 92 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[2]
port 93 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_o[30]
port 94 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 wbs_dat_o[31]
port 95 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[3]
port 96 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[4]
port 97 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[5]
port 98 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_o[6]
port 99 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[7]
port 100 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[8]
port 101 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_o[9]
port 102 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[0]
port 103 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_sel_i[1]
port 104 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_sel_i[2]
port 105 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_sel_i[3]
port 106 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 107 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 108 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 55229 57373
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4136050
string GDS_FILE /mnt/c/Users/Ismael/Efabless-wsl/caravel_tutorial/caravel_example/openlane/SPM_example/runs/SPM_example/results/finishing/SPM_example.magic.gds
string GDS_START 432118
<< end >>

