* NGSPICE file created from SPM_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt SPM_example VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2106_ _2213_/A VGND VGND VPWR VPWR _2194_/A sky130_fd_sc_hd__clkbuf_2
X_2037_ _2285_/A VGND VGND VPWR VPWR _2083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1270_ _1268_/X _1263_/X _1269_/Y VGND VGND VPWR VPWR _1270_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1606_ _2445_/Q _2444_/Q _1606_/C VGND VGND VPWR VPWR _1612_/C sky130_fd_sc_hd__and3_1
X_2586_ _2593_/CLK _2586_/D _2350_/Y VGND VGND VPWR VPWR _2586_/Q sky130_fd_sc_hd__dfrtp_1
X_1537_ input48/X _2429_/Q _1545_/S VGND VGND VPWR VPWR _1538_/A sky130_fd_sc_hd__mux2_1
X_1468_ _1468_/A VGND VGND VPWR VPWR _2469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1399_ _1399_/A VGND VGND VPWR VPWR _2500_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2440_ _2446_/CLK _2440_/D _1923_/Y VGND VGND VPWR VPWR _2440_/Q sky130_fd_sc_hd__dfrtp_1
X_2371_ _2497_/CLK _2371_/D _1837_/Y VGND VGND VPWR VPWR _2371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1322_ _1320_/X _1313_/X _1321_/Y VGND VGND VPWR VPWR _1322_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1253_ input49/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1184_ _1184_/A _1184_/B VGND VGND VPWR VPWR _1187_/B sky130_fd_sc_hd__nor2_1
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2569_ _2575_/CLK _2569_/D _2328_/Y VGND VGND VPWR VPWR _2569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1940_ _1943_/A VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1871_ _1875_/A VGND VGND VPWR VPWR _1871_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2423_ _2561_/CLK _2423_/D _1902_/Y VGND VGND VPWR VPWR _2423_/Q sky130_fd_sc_hd__dfrtp_1
X_2354_ _2354_/A VGND VGND VPWR VPWR _2354_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1305_ _1293_/X _1288_/X _1304_/Y VGND VGND VPWR VPWR _1305_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2285_ _2285_/A _2285_/B _2438_/Q VGND VGND VPWR VPWR _2285_/Y sky130_fd_sc_hd__nor3b_1
X_1236_ _2247_/A VGND VGND VPWR VPWR _2024_/B sky130_fd_sc_hd__buf_2
X_1167_ _1167_/A _1167_/B VGND VGND VPWR VPWR _1168_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _2519_/Q VGND VGND VPWR VPWR _2070_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1923_ _1925_/A VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__inv_2
X_1854_ _1856_/A VGND VGND VPWR VPWR _1854_/Y sky130_fd_sc_hd__inv_2
X_1785_ _2589_/Q _2586_/Q _1784_/B VGND VGND VPWR VPWR _2589_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2406_ _2406_/CLK _2406_/D _1880_/Y VGND VGND VPWR VPWR _2406_/Q sky130_fd_sc_hd__dfrtp_4
X_2337_ _2355_/A VGND VGND VPWR VPWR _2342_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2268_ _2264_/Y _2266_/Y _2267_/X VGND VGND VPWR VPWR _2268_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1219_ _1297_/A VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2199_ _2500_/Q _2198_/X _2165_/X _2189_/X VGND VGND VPWR VPWR _2199_/X sky130_fd_sc_hd__o31a_1
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2497_/CLK sky130_fd_sc_hd__clkbuf_16
X_1570_ input63/X _2414_/Q _1578_/S VGND VGND VPWR VPWR _1571_/A sky130_fd_sc_hd__mux2_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2122_ _2165_/A VGND VGND VPWR VPWR _2122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2053_ _2083_/A _2061_/B _2411_/Q VGND VGND VPWR VPWR _2053_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1906_ _1906_/A VGND VGND VPWR VPWR _1906_/Y sky130_fd_sc_hd__inv_2
X_1837_ _1838_/A VGND VGND VPWR VPWR _1837_/Y sky130_fd_sc_hd__inv_2
X_1768_ _2585_/Q _2582_/Q VGND VGND VPWR VPWR _1768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1699_ _1696_/X _1697_/Y _1706_/C _2414_/Q VGND VGND VPWR VPWR _1700_/B sky130_fd_sc_hd__and4bb_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput75 _2528_/Q VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput97 _2519_/Q VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput86 _2538_/Q VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _1622_/A _1622_/B VGND VGND VPWR VPWR _2370_/D sky130_fd_sc_hd__nor2_1
X_1553_ _1553_/A VGND VGND VPWR VPWR _2422_/D sky130_fd_sc_hd__clkbuf_1
X_1484_ _2461_/Q _2462_/Q _1484_/S VGND VGND VPWR VPWR _1485_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2105_ _2523_/Q VGND VGND VPWR VPWR _2105_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2036_ _2515_/Q VGND VGND VPWR VPWR _2036_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1605_ _1586_/B _1606_/C _1604_/Y VGND VGND VPWR VPWR _2444_/D sky130_fd_sc_hd__a21oi_1
X_2585_ _2589_/CLK _2585_/D _2348_/Y VGND VGND VPWR VPWR _2585_/Q sky130_fd_sc_hd__dfrtp_1
X_1536_ _1558_/A VGND VGND VPWR VPWR _1545_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467_ _2469_/Q _2470_/Q _1473_/S VGND VGND VPWR VPWR _1468_/A sky130_fd_sc_hd__mux2_1
X_1398_ _2500_/Q _2501_/Q _1406_/S VGND VGND VPWR VPWR _1399_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2019_ _2026_/A _2252_/A VGND VGND VPWR VPWR _2231_/A sky130_fd_sc_hd__nand2_2
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _2601_/CLK _2370_/D _1836_/Y VGND VGND VPWR VPWR _2370_/Q sky130_fd_sc_hd__dfrtp_1
X_1321_ _2555_/Q VGND VGND VPWR VPWR _1321_/Y sky130_fd_sc_hd__inv_2
X_1252_ _1374_/A VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1183_ _1183_/A input9/X VGND VGND VPWR VPWR _1187_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2568_ _2568_/CLK _2568_/D _2327_/Y VGND VGND VPWR VPWR _2568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1519_ input56/X _2437_/Q _1523_/S VGND VGND VPWR VPWR _1520_/A sky130_fd_sc_hd__mux2_1
X_2499_ _2503_/CLK _2499_/D _1996_/Y VGND VGND VPWR VPWR _2499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2555_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1870_ _1882_/A VGND VGND VPWR VPWR _1875_/A sky130_fd_sc_hd__buf_2
X_2422_ _2561_/CLK _2422_/D _1900_/Y VGND VGND VPWR VPWR _2422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2353_ _2354_/A VGND VGND VPWR VPWR _2353_/Y sky130_fd_sc_hd__inv_2
X_1304_ _2558_/Q VGND VGND VPWR VPWR _1304_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2284_ _2544_/Q VGND VGND VPWR VPWR _2284_/Y sky130_fd_sc_hd__inv_2
X_1235_ _2026_/A VGND VGND VPWR VPWR _2247_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1166_ _1166_/A _1166_/B VGND VGND VPWR VPWR _1168_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1999_ _1999_/A VGND VGND VPWR VPWR _1999_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1922_ _1925_/A VGND VGND VPWR VPWR _1922_/Y sky130_fd_sc_hd__inv_2
X_1853_ _1856_/A VGND VGND VPWR VPWR _1853_/Y sky130_fd_sc_hd__inv_2
X_1784_ _1784_/A _1784_/B VGND VGND VPWR VPWR _2588_/D sky130_fd_sc_hd__nor2_1
X_2405_ _2587_/CLK _2405_/D _1879_/Y VGND VGND VPWR VPWR _2405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ _2336_/A VGND VGND VPWR VPWR _2336_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2267_ _2508_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2267_/X sky130_fd_sc_hd__o31a_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1218_ _2237_/A VGND VGND VPWR VPWR _1297_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2198_ _2241_/A VGND VGND VPWR VPWR _2198_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2121_ _1673_/C _2118_/X _2119_/X _2120_/Y VGND VGND VPWR VPWR _2121_/Y sky130_fd_sc_hd__o211ai_1
X_2052_ _2517_/Q VGND VGND VPWR VPWR _2052_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1905_ _1906_/A VGND VGND VPWR VPWR _1905_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1836_ _1838_/A VGND VGND VPWR VPWR _1836_/Y sky130_fd_sc_hd__inv_2
X_1767_ _2585_/Q _2582_/Q VGND VGND VPWR VPWR _1767_/X sky130_fd_sc_hd__and2_1
XFILLER_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1698_ _1647_/X _2414_/Q _1696_/X _1697_/Y VGND VGND VPWR VPWR _1700_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2323_/A VGND VGND VPWR VPWR _2319_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput76 _2529_/Q VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput98 _2520_/Q VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput87 _2539_/Q VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1621_ _1643_/A _1621_/B _1621_/C _1621_/D VGND VGND VPWR VPWR _1622_/B sky130_fd_sc_hd__nor4_1
X_1552_ input40/X _2422_/Q _1556_/S VGND VGND VPWR VPWR _1553_/A sky130_fd_sc_hd__mux2_1
X_1483_ _1483_/A VGND VGND VPWR VPWR _2462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2104_ _2097_/Y _2071_/X _2103_/Y VGND VGND VPWR VPWR _2522_/D sky130_fd_sc_hd__o21ai_1
XFILLER_27_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2035_ _2018_/Y _2022_/X _2034_/Y VGND VGND VPWR VPWR _2514_/D sky130_fd_sc_hd__o21ai_1
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1819_ _2601_/Q _2598_/Q VGND VGND VPWR VPWR _1819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1604_ _1586_/B _1606_/C _1194_/X VGND VGND VPWR VPWR _1604_/Y sky130_fd_sc_hd__o21ai_1
X_2584_ _2587_/CLK _2584_/D _2347_/Y VGND VGND VPWR VPWR _2584_/Q sky130_fd_sc_hd__dfrtp_1
X_1535_ _1535_/A VGND VGND VPWR VPWR _2430_/D sky130_fd_sc_hd__clkbuf_1
X_1466_ _1466_/A VGND VGND VPWR VPWR _2470_/D sky130_fd_sc_hd__clkbuf_1
X_1397_ _1430_/A VGND VGND VPWR VPWR _1406_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2018_ _2514_/Q VGND VGND VPWR VPWR _2018_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1320_ _1346_/A VGND VGND VPWR VPWR _1320_/X sky130_fd_sc_hd__clkbuf_2
X_1251_ _1497_/A VGND VGND VPWR VPWR _1374_/A sky130_fd_sc_hd__buf_4
X_1182_ _1182_/A _1182_/B _1182_/C VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__nand3_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_9_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2395_/CLK sky130_fd_sc_hd__clkbuf_16
X_2567_ _2567_/CLK _2567_/D _2326_/Y VGND VGND VPWR VPWR _2567_/Q sky130_fd_sc_hd__dfrtp_1
X_2498_ _2505_/CLK _2498_/D _1995_/Y VGND VGND VPWR VPWR _2498_/Q sky130_fd_sc_hd__dfrtp_1
X_1518_ _1518_/A VGND VGND VPWR VPWR _2438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1449_ _2477_/Q _2478_/Q _1451_/S VGND VGND VPWR VPWR _1450_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2421_ _2561_/CLK _2421_/D _1899_/Y VGND VGND VPWR VPWR _2421_/Q sky130_fd_sc_hd__dfrtp_4
X_2352_ _2354_/A VGND VGND VPWR VPWR _2352_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2283_ _2277_/Y _2246_/X _2282_/Y VGND VGND VPWR VPWR _2543_/D sky130_fd_sc_hd__o21ai_1
X_1303_ input38/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1303_/X sky130_fd_sc_hd__o21ba_1
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1234_ input52/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1234_/X sky130_fd_sc_hd__o21ba_1
XFILLER_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1165_ _1165_/A _1165_/B VGND VGND VPWR VPWR _1165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1998_ _1999_/A VGND VGND VPWR VPWR _1998_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1921_ _1925_/A VGND VGND VPWR VPWR _1921_/Y sky130_fd_sc_hd__inv_2
X_1852_ _1856_/A VGND VGND VPWR VPWR _1852_/Y sky130_fd_sc_hd__inv_2
X_1783_ _1780_/X _1781_/Y _1789_/C _2433_/Q VGND VGND VPWR VPWR _1784_/B sky130_fd_sc_hd__and4bb_1
X_2404_ _2587_/CLK _2404_/D _1878_/Y VGND VGND VPWR VPWR _2404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2335_ _2336_/A VGND VGND VPWR VPWR _2335_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2266_ _1226_/Y _2237_/X _2249_/X _2265_/Y VGND VGND VPWR VPWR _2266_/Y sky130_fd_sc_hd__o211ai_1
X_1217_ _2576_/Q _1209_/X _1211_/X _1216_/Y VGND VGND VPWR VPWR _2575_/D sky130_fd_sc_hd__a22o_1
X_2197_ _1269_/Y _2135_/X _2162_/X _2196_/Y VGND VGND VPWR VPWR _2197_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2120_ _2144_/A _2459_/Q VGND VGND VPWR VPWR _2120_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2503_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2051_ _2045_/Y _2022_/X _2050_/Y VGND VGND VPWR VPWR _2516_/D sky130_fd_sc_hd__o21ai_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1904_ _1906_/A VGND VGND VPWR VPWR _1904_/Y sky130_fd_sc_hd__inv_2
X_1835_ _1838_/A VGND VGND VPWR VPWR _1835_/Y sky130_fd_sc_hd__inv_2
X_1766_ _2583_/Q _2580_/Q _1765_/B VGND VGND VPWR VPWR _2583_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1697_ _2393_/Q _2390_/Q VGND VGND VPWR VPWR _1697_/Y sky130_fd_sc_hd__nor2_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2324_/A VGND VGND VPWR VPWR _2323_/A sky130_fd_sc_hd__buf_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2249_ _2249_/A VGND VGND VPWR VPWR _2249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput99 _2521_/Q VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput77 _2530_/Q VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput88 _2540_/Q VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1620_ _1828_/A _1621_/C _1621_/D _1621_/B VGND VGND VPWR VPWR _1622_/A sky130_fd_sc_hd__o22a_1
X_1551_ _1551_/A VGND VGND VPWR VPWR _2423_/D sky130_fd_sc_hd__clkbuf_1
X_1482_ _2462_/Q _2463_/Q _1484_/S VGND VGND VPWR VPWR _1483_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2103_ _2098_/Y _2100_/Y _2102_/X VGND VGND VPWR VPWR _2103_/Y sky130_fd_sc_hd__o21ai_2
X_2034_ _2024_/Y _2031_/Y _2033_/Y VGND VGND VPWR VPWR _2034_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_35_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1818_ _2601_/Q _2598_/Q VGND VGND VPWR VPWR _1818_/X sky130_fd_sc_hd__and2_1
XFILLER_2_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1749_ _2579_/Q _2404_/Q VGND VGND VPWR VPWR _1749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1603_ _1603_/A VGND VGND VPWR VPWR _2443_/D sky130_fd_sc_hd__clkbuf_1
X_2583_ _2589_/CLK _2583_/D _2346_/Y VGND VGND VPWR VPWR _2583_/Q sky130_fd_sc_hd__dfrtp_1
X_1534_ input49/X _2430_/Q _1534_/S VGND VGND VPWR VPWR _1535_/A sky130_fd_sc_hd__mux2_1
X_1465_ _2470_/Q _2471_/Q _1473_/S VGND VGND VPWR VPWR _1466_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ _1396_/A VGND VGND VPWR VPWR _2501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ _1214_/X _2016_/X _2513_/Q VGND VGND VPWR VPWR _2513_/D sky130_fd_sc_hd__a21oi_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1250_ _2570_/Q _1233_/X _1247_/X _1249_/Y VGND VGND VPWR VPWR _2569_/D sky130_fd_sc_hd__a22o_1
X_1181_ input4/X input3/X VGND VGND VPWR VPWR _1182_/C sky130_fd_sc_hd__nor2_1
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2566_ _2567_/CLK _2566_/D _2325_/Y VGND VGND VPWR VPWR _2566_/Q sky130_fd_sc_hd__dfrtp_1
X_1517_ input58/X _2438_/Q _1523_/S VGND VGND VPWR VPWR _1518_/A sky130_fd_sc_hd__mux2_1
X_2497_ _2497_/CLK _2497_/D _1993_/Y VGND VGND VPWR VPWR _2497_/Q sky130_fd_sc_hd__dfrtp_1
X_1448_ _1448_/A VGND VGND VPWR VPWR _2478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1379_ _2508_/Q _2509_/Q _1383_/S VGND VGND VPWR VPWR _1380_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ _2560_/CLK _2420_/D _1898_/Y VGND VGND VPWR VPWR _2420_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2351_ _2354_/A VGND VGND VPWR VPWR _2351_/Y sky130_fd_sc_hd__inv_2
X_1302_ _1374_/A VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__clkbuf_1
X_2282_ _2278_/Y _2280_/Y _2281_/X VGND VGND VPWR VPWR _2282_/Y sky130_fd_sc_hd__o21ai_2
X_1233_ _1608_/B VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1164_ _1200_/A VGND VGND VPWR VPWR _2213_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1997_ _1999_/A VGND VGND VPWR VPWR _1997_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2549_ _2549_/CLK _2549_/D _2304_/Y VGND VGND VPWR VPWR _2549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1920_ _1944_/A VGND VGND VPWR VPWR _1925_/A sky130_fd_sc_hd__buf_4
X_1851_ _2367_/A VGND VGND VPWR VPWR _1856_/A sky130_fd_sc_hd__buf_2
X_1782_ _1747_/X _2433_/Q _1780_/X _1781_/Y VGND VGND VPWR VPWR _1784_/A sky130_fd_sc_hd__o2bb2a_1
X_2403_ _2403_/CLK _2403_/D _1877_/Y VGND VGND VPWR VPWR _2403_/Q sky130_fd_sc_hd__dfrtp_1
X_2334_ _2336_/A VGND VGND VPWR VPWR _2334_/Y sky130_fd_sc_hd__inv_2
X_2265_ _2272_/A _2476_/Q VGND VGND VPWR VPWR _2265_/Y sky130_fd_sc_hd__nand2_1
X_1216_ _1212_/X _1214_/X _1215_/Y VGND VGND VPWR VPWR _1216_/Y sky130_fd_sc_hd__o21ai_1
X_2196_ _2229_/A _2468_/Q VGND VGND VPWR VPWR _2196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2050_ _2046_/Y _2048_/Y _2049_/X VGND VGND VPWR VPWR _2050_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _1906_/A VGND VGND VPWR VPWR _1903_/Y sky130_fd_sc_hd__inv_2
X_1834_ _1838_/A VGND VGND VPWR VPWR _1834_/Y sky130_fd_sc_hd__inv_2
X_1765_ _1765_/A _1765_/B VGND VGND VPWR VPWR _2582_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1696_ _2393_/Q _2390_/Q VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__and2_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2317_/A VGND VGND VPWR VPWR _2317_/Y sky130_fd_sc_hd__inv_2
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2264_/A _2285_/B _2433_/Q VGND VGND VPWR VPWR _2248_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2179_ _2187_/A _2466_/Q VGND VGND VPWR VPWR _2179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput78 _2531_/Q VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput89 _2541_/Q VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1550_ input41/X _2423_/Q _1556_/S VGND VGND VPWR VPWR _1551_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1481_ _1481_/A VGND VGND VPWR VPWR _2463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2102_ _2489_/Q _2066_/X _2078_/X _2101_/X VGND VGND VPWR VPWR _2102_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2033_ _2481_/Q _2074_/A _2032_/X VGND VGND VPWR VPWR _2033_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1817_ _2599_/Q _2596_/Q _1816_/B VGND VGND VPWR VPWR _2599_/D sky130_fd_sc_hd__a21o_1
X_1748_ _2579_/Q _2404_/Q VGND VGND VPWR VPWR _1748_/X sky130_fd_sc_hd__and2_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1679_ _1676_/X _1677_/Y _1706_/C _2417_/Q VGND VGND VPWR VPWR _1680_/B sky130_fd_sc_hd__and4bb_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1602_ _1606_/C _1614_/C _1602_/C VGND VGND VPWR VPWR _1603_/A sky130_fd_sc_hd__and3b_1
X_2582_ _2589_/CLK _2582_/D _2345_/Y VGND VGND VPWR VPWR _2582_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1533_ _1533_/A VGND VGND VPWR VPWR _2431_/D sky130_fd_sc_hd__clkbuf_1
X_1464_ _1486_/A VGND VGND VPWR VPWR _1473_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1395_ _2501_/Q _2502_/Q _1395_/S VGND VGND VPWR VPWR _1396_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2016_ _2252_/A VGND VGND VPWR VPWR _2016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1182_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2565_ _2567_/CLK _2565_/D _2323_/Y VGND VGND VPWR VPWR _2565_/Q sky130_fd_sc_hd__dfrtp_1
X_1516_ _1516_/A VGND VGND VPWR VPWR _2439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2496_ _2496_/CLK _2496_/D _1992_/Y VGND VGND VPWR VPWR _2496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1447_ _2478_/Q _2479_/Q _1451_/S VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__mux2_1
X_1378_ _1378_/A VGND VGND VPWR VPWR _2509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _2354_/A VGND VGND VPWR VPWR _2350_/Y sky130_fd_sc_hd__inv_2
X_1301_ _2560_/Q _1286_/X _1298_/X _1300_/Y VGND VGND VPWR VPWR _2559_/D sky130_fd_sc_hd__a22o_1
X_2281_ _2510_/Q _2066_/A _2252_/X _2032_/X VGND VGND VPWR VPWR _2281_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1232_ _2573_/Q _1209_/X _1229_/X _1231_/Y VGND VGND VPWR VPWR _2572_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1996_ _1999_/A VGND VGND VPWR VPWR _1996_/Y sky130_fd_sc_hd__inv_2
X_2548_ _2550_/CLK _2548_/D _2303_/Y VGND VGND VPWR VPWR _2548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2479_ _2504_/CLK _2479_/D _1971_/Y VGND VGND VPWR VPWR _2479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1850_ _1850_/A VGND VGND VPWR VPWR _1850_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1781_ _2589_/Q _2586_/Q VGND VGND VPWR VPWR _1781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2402_ _2487_/CLK _2402_/D _1875_/Y VGND VGND VPWR VPWR _2402_/Q sky130_fd_sc_hd__dfrtp_1
X_2333_ _2336_/A VGND VGND VPWR VPWR _2333_/Y sky130_fd_sc_hd__inv_2
X_2264_ _2264_/A _2285_/B _2435_/Q VGND VGND VPWR VPWR _2264_/Y sky130_fd_sc_hd__nor3b_1
X_1215_ _2575_/Q VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__inv_2
X_2195_ _2238_/A VGND VGND VPWR VPWR _2229_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1979_ _1980_/A VGND VGND VPWR VPWR _1979_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _1906_/A VGND VGND VPWR VPWR _1902_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2529_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1833_ _2367_/A VGND VGND VPWR VPWR _1838_/A sky130_fd_sc_hd__buf_2
X_1764_ _1761_/X _1762_/Y _1789_/C _2436_/Q VGND VGND VPWR VPWR _1765_/B sky130_fd_sc_hd__and4bb_1
X_1695_ _2391_/Q _2388_/Q _1694_/B VGND VGND VPWR VPWR _2391_/D sky130_fd_sc_hd__a21o_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2317_/A VGND VGND VPWR VPWR _2316_/Y sky130_fd_sc_hd__inv_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2247_/A VGND VGND VPWR VPWR _2285_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2178_ _2178_/A _2228_/B VGND VGND VPWR VPWR _2178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput79 _2532_/Q VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1480_ _2463_/Q _2464_/Q _1484_/S VGND VGND VPWR VPWR _1481_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2101_ _2146_/A VGND VGND VPWR VPWR _2101_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2032_ _2231_/A VGND VGND VPWR VPWR _2032_/X sky130_fd_sc_hd__buf_2
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1816_ _1816_/A _1816_/B VGND VGND VPWR VPWR _2598_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1747_ _1747_/A VGND VGND VPWR VPWR _1747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1678_ _1647_/X _2417_/Q _1676_/X _1677_/Y VGND VGND VPWR VPWR _1680_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1601_ _1588_/A _1593_/A _2442_/Q _2443_/Q VGND VGND VPWR VPWR _1602_/C sky130_fd_sc_hd__a31o_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2581_ _2587_/CLK _2581_/D _2344_/Y VGND VGND VPWR VPWR _2581_/Q sky130_fd_sc_hd__dfrtp_1
X_1532_ input50/X _2431_/Q _1534_/S VGND VGND VPWR VPWR _1533_/A sky130_fd_sc_hd__mux2_1
X_1463_ _1463_/A VGND VGND VPWR VPWR _2471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1394_ _1394_/A VGND VGND VPWR VPWR _2502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2015_ _2028_/B _2028_/C _2028_/D VGND VGND VPWR VPWR _2252_/A sky130_fd_sc_hd__nand3_4
XFILLER_50_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2564_ _2567_/CLK _2564_/D _2322_/Y VGND VGND VPWR VPWR _2564_/Q sky130_fd_sc_hd__dfrtp_1
X_1515_ input59/X _2439_/Q _1523_/S VGND VGND VPWR VPWR _1516_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2495_ _2495_/CLK _2495_/D _1991_/Y VGND VGND VPWR VPWR _2495_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1446_ _1446_/A VGND VGND VPWR VPWR _2479_/D sky130_fd_sc_hd__clkbuf_1
X_1377_ _2509_/Q _2510_/Q _1383_/S VGND VGND VPWR VPWR _1378_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1300_ _1293_/X _1288_/X _1299_/Y VGND VGND VPWR VPWR _1300_/Y sky130_fd_sc_hd__o21ai_1
X_2280_ _1215_/Y _2237_/X _2249_/X _2279_/Y VGND VGND VPWR VPWR _2280_/Y sky130_fd_sc_hd__o211ai_1
X_1231_ _1212_/X _1214_/X _2257_/A VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _1999_/A VGND VGND VPWR VPWR _1995_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2547_ _2550_/CLK _2547_/D _2302_/Y VGND VGND VPWR VPWR _2547_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2478_ _2504_/CLK _2478_/D _1970_/Y VGND VGND VPWR VPWR _2478_/Q sky130_fd_sc_hd__dfrtp_1
X_1429_ _1429_/A VGND VGND VPWR VPWR _2486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1780_ _2589_/Q _2586_/Q VGND VGND VPWR VPWR _1780_/X sky130_fd_sc_hd__and2_1
X_2401_ _2403_/CLK _2401_/D _1874_/Y VGND VGND VPWR VPWR _2401_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2332_ _2336_/A VGND VGND VPWR VPWR _2332_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2263_ _2541_/Q VGND VGND VPWR VPWR _2263_/Y sky130_fd_sc_hd__inv_2
X_1214_ _2054_/A VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__buf_4
X_2194_ _2194_/A _2236_/B _2427_/Q VGND VGND VPWR VPWR _2194_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1978_ _1980_/A VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_2_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _1913_/A VGND VGND VPWR VPWR _1906_/A sky130_fd_sc_hd__buf_2
X_1832_ _2361_/A VGND VGND VPWR VPWR _2367_/A sky130_fd_sc_hd__clkbuf_2
X_1763_ _1747_/X _2436_/Q _1761_/X _1762_/Y VGND VGND VPWR VPWR _1765_/A sky130_fd_sc_hd__o2bb2a_1
X_1694_ _1694_/A _1694_/B VGND VGND VPWR VPWR _2390_/D sky130_fd_sc_hd__nor2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2317_/A VGND VGND VPWR VPWR _2315_/Y sky130_fd_sc_hd__inv_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2246_/A VGND VGND VPWR VPWR _2246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2177_ _2531_/Q VGND VGND VPWR VPWR _2177_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput69 _2513_/Q VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2100_ _1686_/C _1583_/S _2074_/X _2099_/Y VGND VGND VPWR VPWR _2100_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2031_ _1672_/A _2292_/B _2027_/Y _2030_/X VGND VGND VPWR VPWR _2031_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ _1828_/A _1815_/B _1815_/C _1815_/D VGND VGND VPWR VPWR _1816_/B sky130_fd_sc_hd__nor4_1
X_1746_ _2407_/Q _2402_/Q _1745_/B VGND VGND VPWR VPWR _2407_/D sky130_fd_sc_hd__a21o_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1677_ _2387_/Q _2384_/Q VGND VGND VPWR VPWR _1677_/Y sky130_fd_sc_hd__nor2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _2229_/A _2472_/Q VGND VGND VPWR VPWR _2229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1600_ _2441_/Q _2440_/Q _2443_/Q _2442_/Q VGND VGND VPWR VPWR _1606_/C sky130_fd_sc_hd__and4_1
X_2580_ _2587_/CLK _2580_/D _2342_/Y VGND VGND VPWR VPWR _2580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1531_ _1531_/A VGND VGND VPWR VPWR _2432_/D sky130_fd_sc_hd__clkbuf_1
X_1462_ _2471_/Q _2472_/Q _1462_/S VGND VGND VPWR VPWR _1463_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1393_ _2502_/Q _2503_/Q _1395_/S VGND VGND VPWR VPWR _1394_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2014_ _2014_/A _2014_/B VGND VGND VPWR VPWR _2028_/D sky130_fd_sc_hd__nor2_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1729_ _2401_/Q _2398_/Q _1728_/B VGND VGND VPWR VPWR _2401_/D sky130_fd_sc_hd__a21o_1
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2563_ _2567_/CLK _2563_/D _2321_/Y VGND VGND VPWR VPWR _2563_/Q sky130_fd_sc_hd__dfrtp_1
X_1514_ _1558_/A VGND VGND VPWR VPWR _1523_/S sky130_fd_sc_hd__buf_2
X_2494_ _2496_/CLK _2494_/D _1990_/Y VGND VGND VPWR VPWR _2494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1445_ _2479_/Q _2480_/Q _1451_/S VGND VGND VPWR VPWR _1446_/A sky130_fd_sc_hd__mux2_1
X_1376_ _1376_/A VGND VGND VPWR VPWR _2510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _2572_/Q VGND VGND VPWR VPWR _2257_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ _2006_/A VGND VGND VPWR VPWR _1999_/A sky130_fd_sc_hd__buf_2
X_2546_ _2553_/CLK _2546_/D _2301_/Y VGND VGND VPWR VPWR _2546_/Q sky130_fd_sc_hd__dfrtp_4
X_2477_ _2587_/CLK _2477_/D _1968_/Y VGND VGND VPWR VPWR _2477_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1428_ _2486_/Q _2487_/Q _1428_/S VGND VGND VPWR VPWR _1429_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1359_ _2549_/Q _1339_/X _1356_/X _1358_/Y VGND VGND VPWR VPWR _2548_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2400_ _2403_/CLK _2400_/D _1873_/Y VGND VGND VPWR VPWR _2400_/Q sky130_fd_sc_hd__dfrtp_1
X_2331_ _2355_/A VGND VGND VPWR VPWR _2336_/A sky130_fd_sc_hd__buf_2
X_2262_ _2256_/Y _2246_/X _2261_/Y VGND VGND VPWR VPWR _2540_/D sky130_fd_sc_hd__o21ai_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1213_ _2238_/A VGND VGND VPWR VPWR _2054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2193_ _2533_/Q VGND VGND VPWR VPWR _2193_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ _1980_/A VGND VGND VPWR VPWR _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2529_ _2529_/CLK _2529_/D VGND VGND VPWR VPWR _2529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ _1900_/A VGND VGND VPWR VPWR _1900_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ input1/X VGND VGND VPWR VPWR _2361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1762_ _2583_/Q _2580_/Q VGND VGND VPWR VPWR _1762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1693_ _1777_/A _1693_/B _1693_/C _1693_/D VGND VGND VPWR VPWR _1694_/B sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2549_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2314_ _2317_/A VGND VGND VPWR VPWR _2314_/Y sky130_fd_sc_hd__inv_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _2539_/Q VGND VGND VPWR VPWR _2245_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2176_ _2169_/Y _2160_/X _2175_/Y VGND VGND VPWR VPWR _2530_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ _2074_/A VGND VGND VPWR VPWR _2030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1814_ _1722_/X _1815_/C _1815_/D _1815_/B VGND VGND VPWR VPWR _1816_/A sky130_fd_sc_hd__o22a_1
X_1745_ _1745_/A _1745_/B VGND VGND VPWR VPWR _2406_/D sky130_fd_sc_hd__nor2_1
X_1676_ _2387_/Q _2384_/Q VGND VGND VPWR VPWR _1676_/X sky130_fd_sc_hd__and2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2228_ _2228_/A _2228_/B VGND VGND VPWR VPWR _2228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2159_ _2529_/Q VGND VGND VPWR VPWR _2159_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1530_ input51/X _2432_/Q _1534_/S VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__mux2_1
X_1461_ _1461_/A VGND VGND VPWR VPWR _2472_/D sky130_fd_sc_hd__clkbuf_1
X_1392_ _1392_/A VGND VGND VPWR VPWR _2503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2013_ _2013_/A _2013_/B VGND VGND VPWR VPWR _2014_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1728_ _1728_/A _1728_/B VGND VGND VPWR VPWR _2400_/D sky130_fd_sc_hd__nor2_1
X_1659_ _1655_/X _1656_/Y _1706_/C _2420_/Q VGND VGND VPWR VPWR _1660_/B sky130_fd_sc_hd__and4bb_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2562_ _2567_/CLK _2562_/D _2320_/Y VGND VGND VPWR VPWR _2562_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1513_ _2186_/A VGND VGND VPWR VPWR _1558_/A sky130_fd_sc_hd__buf_2
X_2493_ _2495_/CLK _2493_/D _1989_/Y VGND VGND VPWR VPWR _2493_/Q sky130_fd_sc_hd__dfrtp_1
X_1444_ _1444_/A VGND VGND VPWR VPWR _2480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1375_ _2510_/Q _2511_/Q _1383_/S VGND VGND VPWR VPWR _1376_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1993_ _1993_/A VGND VGND VPWR VPWR _1993_/Y sky130_fd_sc_hd__inv_2
X_2545_ _2573_/CLK _2545_/D VGND VGND VPWR VPWR _2545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2476_ _2578_/CLK _2476_/D _1967_/Y VGND VGND VPWR VPWR _2476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1427_ _1427_/A VGND VGND VPWR VPWR _2487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1358_ _1346_/X _1341_/X _2046_/A VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1289_ _2561_/Q VGND VGND VPWR VPWR _2161_/A sky130_fd_sc_hd__inv_2
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2330_ input1/X VGND VGND VPWR VPWR _2355_/A sky130_fd_sc_hd__buf_4
X_2261_ _2257_/Y _2259_/Y _2260_/X VGND VGND VPWR VPWR _2261_/Y sky130_fd_sc_hd__o21ai_2
X_1212_ _1293_/A VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__clkbuf_2
X_2192_ _2184_/Y _2160_/X _2191_/Y VGND VGND VPWR VPWR _2532_/D sky130_fd_sc_hd__o21ai_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1976_ _1980_/A VGND VGND VPWR VPWR _1976_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2528_ _2528_/CLK _2528_/D VGND VGND VPWR VPWR _2528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2459_ _2487_/CLK _2459_/D _1946_/Y VGND VGND VPWR VPWR _2459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ _2369_/Q _2600_/Q _1829_/B VGND VGND VPWR VPWR _2369_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1761_ _2583_/Q _2580_/Q VGND VGND VPWR VPWR _1761_/X sky130_fd_sc_hd__and2_1
X_1692_ _1631_/X _1693_/C _1693_/D _1693_/B VGND VGND VPWR VPWR _1694_/A sky130_fd_sc_hd__o22a_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2317_/A VGND VGND VPWR VPWR _2313_/Y sky130_fd_sc_hd__inv_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2235_/Y _2203_/X _2243_/Y VGND VGND VPWR VPWR _2538_/D sky130_fd_sc_hd__o21ai_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2387_/CLK sky130_fd_sc_hd__clkbuf_16
X_2175_ _2171_/Y _2173_/Y _2174_/X VGND VGND VPWR VPWR _2175_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1959_ _1962_/A VGND VGND VPWR VPWR _1959_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1813_ _2599_/Q _2596_/Q VGND VGND VPWR VPWR _1815_/B sky130_fd_sc_hd__nor2_1
X_1744_ _1741_/X _1742_/Y _1751_/C _2408_/Q VGND VGND VPWR VPWR _1745_/B sky130_fd_sc_hd__and4bb_1
X_1675_ _2385_/Q _2382_/Q _1674_/B VGND VGND VPWR VPWR _2385_/D sky130_fd_sc_hd__a21o_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2537_/Q VGND VGND VPWR VPWR _2227_/Y sky130_fd_sc_hd__inv_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2158_ _2150_/Y _2116_/X _2157_/Y VGND VGND VPWR VPWR _2528_/D sky130_fd_sc_hd__o21ai_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2089_ _2521_/Q VGND VGND VPWR VPWR _2089_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1460_ _2472_/Q _2473_/Q _1462_/S VGND VGND VPWR VPWR _1461_/A sky130_fd_sc_hd__mux2_1
X_1391_ _2503_/Q _2504_/Q _1395_/S VGND VGND VPWR VPWR _1392_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2012_ _2448_/Q _2012_/B VGND VGND VPWR VPWR _2013_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1727_ _1777_/A _1727_/B _1727_/C _1727_/D VGND VGND VPWR VPWR _1728_/B sky130_fd_sc_hd__nor4_1
X_1658_ _1747_/A VGND VGND VPWR VPWR _1706_/C sky130_fd_sc_hd__clkbuf_2
X_1589_ _1589_/A VGND VGND VPWR VPWR _1614_/C sky130_fd_sc_hd__clkbuf_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2561_ _2561_/CLK _2561_/D _2319_/Y VGND VGND VPWR VPWR _2561_/Q sky130_fd_sc_hd__dfrtp_1
X_1512_ _1512_/A _2028_/B _2028_/C _1512_/D VGND VGND VPWR VPWR _2186_/A sky130_fd_sc_hd__nand4_4
X_2492_ _2492_/CLK _2492_/D _1987_/Y VGND VGND VPWR VPWR _2492_/Q sky130_fd_sc_hd__dfrtp_1
X_1443_ _2480_/Q _2481_/Q _1451_/S VGND VGND VPWR VPWR _1444_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1374_ _1374_/A VGND VGND VPWR VPWR _1383_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1992_ _1993_/A VGND VGND VPWR VPWR _1992_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2560_/CLK sky130_fd_sc_hd__clkbuf_16
X_2544_ _2573_/CLK _2544_/D VGND VGND VPWR VPWR _2544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2475_ _2578_/CLK _2475_/D _1966_/Y VGND VGND VPWR VPWR _2475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1426_ _2487_/Q _2488_/Q _1428_/S VGND VGND VPWR VPWR _1427_/A sky130_fd_sc_hd__mux2_1
X_1357_ _2548_/Q VGND VGND VPWR VPWR _2046_/A sky130_fd_sc_hd__inv_2
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1288_ _2024_/B VGND VGND VPWR VPWR _1288_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2260_ _2507_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2260_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1211_ input56/X _1191_/X _1339_/A VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__o21ba_1
X_2191_ _2185_/Y _2188_/Y _2190_/X VGND VGND VPWR VPWR _2191_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ _1975_/A VGND VGND VPWR VPWR _1980_/A sky130_fd_sc_hd__buf_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2527_ _2528_/CLK _2527_/D VGND VGND VPWR VPWR _2527_/Q sky130_fd_sc_hd__dfxtp_1
X_2458_ _2487_/CLK _2458_/D _1945_/Y VGND VGND VPWR VPWR _2458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1409_ _2495_/Q _2496_/Q _1417_/S VGND VGND VPWR VPWR _1410_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2389_ _2395_/CLK _2389_/D _1860_/Y VGND VGND VPWR VPWR _2389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1760_ _2581_/Q _2578_/Q _1759_/B VGND VGND VPWR VPWR _2581_/D sky130_fd_sc_hd__a21o_1
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1691_ _2391_/Q _2388_/Q VGND VGND VPWR VPWR _1693_/B sky130_fd_sc_hd__nor2_1
X_2312_ _2324_/A VGND VGND VPWR VPWR _2317_/A sky130_fd_sc_hd__buf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2243_ _2236_/Y _2240_/Y _2242_/X VGND VGND VPWR VPWR _2243_/Y sky130_fd_sc_hd__o21ai_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _2497_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2174_/X sky130_fd_sc_hd__o31a_1
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1958_ _1962_/A VGND VGND VPWR VPWR _1958_/Y sky130_fd_sc_hd__inv_2
X_1889_ _1913_/A VGND VGND VPWR VPWR _1894_/A sky130_fd_sc_hd__buf_2
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_79_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1812_ _2599_/Q _2596_/Q VGND VGND VPWR VPWR _1815_/D sky130_fd_sc_hd__and2_1
X_1743_ _1702_/X _2408_/Q _1741_/X _1742_/Y VGND VGND VPWR VPWR _1745_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1674_ _1674_/A _1674_/B VGND VGND VPWR VPWR _2384_/D sky130_fd_sc_hd__nor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2220_/Y _2203_/X _2225_/Y VGND VGND VPWR VPWR _2536_/D sky130_fd_sc_hd__o21ai_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2157_ _2151_/Y _2154_/Y _2156_/X VGND VGND VPWR VPWR _2157_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2088_ _2082_/Y _2071_/X _2087_/Y VGND VGND VPWR VPWR _2520_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1390_ _1390_/A VGND VGND VPWR VPWR _2504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2011_ _2011_/A VGND VGND VPWR VPWR _2011_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1726_ _1722_/X _1727_/C _1727_/D _1727_/B VGND VGND VPWR VPWR _1728_/A sky130_fd_sc_hd__o22a_1
X_1657_ _1647_/X _2420_/Q _1655_/X _1656_/Y VGND VGND VPWR VPWR _1660_/A sky130_fd_sc_hd__o2bb2a_1
X_1588_ _1588_/A _2440_/Q _2443_/Q _2442_/Q VGND VGND VPWR VPWR _1588_/X sky130_fd_sc_hd__or4_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2209_ _2501_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2209_/X sky130_fd_sc_hd__o31a_1
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2560_ _2560_/CLK _2560_/D _2317_/Y VGND VGND VPWR VPWR _2560_/Q sky130_fd_sc_hd__dfrtp_1
X_2491_ _2495_/CLK _2491_/D _1986_/Y VGND VGND VPWR VPWR _2491_/Q sky130_fd_sc_hd__dfrtp_1
X_1511_ _1511_/A VGND VGND VPWR VPWR _2449_/D sky130_fd_sc_hd__clkbuf_1
X_1442_ _1486_/A VGND VGND VPWR VPWR _1451_/S sky130_fd_sc_hd__clkbuf_2
X_1373_ _1373_/A VGND VGND VPWR VPWR _2511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1709_ _2397_/Q _2394_/Q VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__and2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1991_ _1993_/A VGND VGND VPWR VPWR _1991_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2543_ _2573_/CLK _2543_/D VGND VGND VPWR VPWR _2543_/Q sky130_fd_sc_hd__dfxtp_1
X_2474_ _2504_/CLK _2474_/D _1965_/Y VGND VGND VPWR VPWR _2474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ _1425_/A VGND VGND VPWR VPWR _2488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1356_ input57/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1356_/X sky130_fd_sc_hd__o21ba_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1287_ input41/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__o21ba_1
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1210_ _1199_/Y _1207_/X _1209_/X _2577_/Q VGND VGND VPWR VPWR _2576_/D sky130_fd_sc_hd__a2bb2o_1
X_2190_ _2499_/Q _2155_/X _2165_/X _2189_/X VGND VGND VPWR VPWR _2190_/X sky130_fd_sc_hd__o31a_1
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1974_ _1974_/A VGND VGND VPWR VPWR _1974_/Y sky130_fd_sc_hd__inv_2
X_2526_ _2528_/CLK _2526_/D VGND VGND VPWR VPWR _2526_/Q sky130_fd_sc_hd__dfxtp_1
X_2457_ _2484_/CLK _2457_/D _1943_/Y VGND VGND VPWR VPWR _2457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1408_ _1430_/A VGND VGND VPWR VPWR _1417_/S sky130_fd_sc_hd__clkbuf_2
X_2388_ _2406_/CLK _2388_/D _1859_/Y VGND VGND VPWR VPWR _2388_/Q sky130_fd_sc_hd__dfrtp_1
X_1339_ _1339_/A VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1690_ _2391_/Q _2388_/Q VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__and2_1
X_2311_ _2311_/A VGND VGND VPWR VPWR _2311_/Y sky130_fd_sc_hd__inv_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2242_ _2505_/Q _2241_/X _2208_/X _2231_/X VGND VGND VPWR VPWR _2242_/X sky130_fd_sc_hd__o31a_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2173_ _1628_/C _2118_/X _2162_/X _2172_/Y VGND VGND VPWR VPWR _2173_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_65_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1957_ _1975_/A VGND VGND VPWR VPWR _1962_/A sky130_fd_sc_hd__buf_2
X_1888_ _2361_/A VGND VGND VPWR VPWR _1913_/A sky130_fd_sc_hd__clkbuf_4
X_2509_ _2510_/CLK _2509_/D _2008_/Y VGND VGND VPWR VPWR _2509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ _2428_/Q VGND VGND VPWR VPWR _1815_/C sky130_fd_sc_hd__clkinv_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1742_ _2407_/Q _2402_/Q VGND VGND VPWR VPWR _1742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1673_ _1777_/A _1673_/B _1673_/C _1673_/D VGND VGND VPWR VPWR _1674_/B sky130_fd_sc_hd__nor4_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2221_/Y _2223_/Y _2224_/X VGND VGND VPWR VPWR _2225_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2156_ _2495_/Q _2155_/X _2122_/X _2146_/X VGND VGND VPWR VPWR _2156_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2087_ _2083_/Y _2085_/Y _2086_/X VGND VGND VPWR VPWR _2087_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2010_ _2011_/A VGND VGND VPWR VPWR _2010_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1725_ _2401_/Q _2398_/Q VGND VGND VPWR VPWR _1727_/B sky130_fd_sc_hd__nor2_1
X_1656_ _2381_/Q _2378_/Q VGND VGND VPWR VPWR _1656_/Y sky130_fd_sc_hd__nor2_1
X_1587_ _2441_/Q VGND VGND VPWR VPWR _1588_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2252_/A VGND VGND VPWR VPWR _2208_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2139_ _2134_/Y _2137_/Y _2138_/X VGND VGND VPWR VPWR _2139_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2490_ _2492_/CLK _2490_/D _1985_/Y VGND VGND VPWR VPWR _2490_/Q sky130_fd_sc_hd__dfrtp_1
X_1510_ _2449_/Q _2450_/Q _1589_/A VGND VGND VPWR VPWR _1511_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1441_ _2448_/Q VGND VGND VPWR VPWR _1486_/A sky130_fd_sc_hd__buf_2
X_1372_ _2511_/Q _2512_/Q _1372_/S VGND VGND VPWR VPWR _1373_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1708_ _2395_/Q _2392_/Q _1707_/B VGND VGND VPWR VPWR _2395_/D sky130_fd_sc_hd__a21o_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1639_ _2422_/Q VGND VGND VPWR VPWR _1643_/C sky130_fd_sc_hd__clkinv_2
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1990_ _1993_/A VGND VGND VPWR VPWR _1990_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2542_ _2573_/CLK _2542_/D VGND VGND VPWR VPWR _2542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2473_ _2504_/CLK _2473_/D _1964_/Y VGND VGND VPWR VPWR _2473_/Q sky130_fd_sc_hd__dfrtp_1
X_1424_ _2488_/Q _2489_/Q _1428_/S VGND VGND VPWR VPWR _1425_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1355_ _1497_/A VGND VGND VPWR VPWR _1372_/S sky130_fd_sc_hd__buf_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1608_/B VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1973_ _1974_/A VGND VGND VPWR VPWR _1973_/Y sky130_fd_sc_hd__inv_2
X_2525_ _2528_/CLK _2525_/D VGND VGND VPWR VPWR _2525_/Q sky130_fd_sc_hd__dfxtp_1
X_2456_ _2484_/CLK _2456_/D _1942_/Y VGND VGND VPWR VPWR _2456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1407_ _1407_/A VGND VGND VPWR VPWR _2496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2387_ _2387_/CLK _2387_/D _1856_/Y VGND VGND VPWR VPWR _2387_/Q sky130_fd_sc_hd__dfrtp_1
X_1338_ _2553_/Q _1311_/X _1335_/X _1337_/Y VGND VGND VPWR VPWR _2552_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1269_ _2565_/Q VGND VGND VPWR VPWR _1269_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2310_ _2311_/A VGND VGND VPWR VPWR _2310_/Y sky130_fd_sc_hd__inv_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2241_/A VGND VGND VPWR VPWR _2241_/X sky130_fd_sc_hd__clkbuf_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2172_ _2187_/A _2465_/Q VGND VGND VPWR VPWR _2172_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1956_ _1956_/A VGND VGND VPWR VPWR _1956_/Y sky130_fd_sc_hd__inv_2
X_1887_ _1887_/A VGND VGND VPWR VPWR _1887_/Y sky130_fd_sc_hd__inv_2
X_2508_ _2510_/CLK _2508_/D _2007_/Y VGND VGND VPWR VPWR _2508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2439_ _2578_/CLK _2439_/D _1922_/Y VGND VGND VPWR VPWR _2439_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ _2597_/Q _2594_/Q _1809_/B VGND VGND VPWR VPWR _2597_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1741_ _2407_/Q _2402_/Q VGND VGND VPWR VPWR _1741_/X sky130_fd_sc_hd__and2_1
XFILLER_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1672_ _1672_/A VGND VGND VPWR VPWR _1777_/A sky130_fd_sc_hd__clkbuf_4
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2503_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2224_/X sky130_fd_sc_hd__o31a_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2155_ _2241_/A VGND VGND VPWR VPWR _2155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2086_ _2487_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2086_/X sky130_fd_sc_hd__o31a_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1939_ _1943_/A VGND VGND VPWR VPWR _1939_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1724_ _2401_/Q _2398_/Q VGND VGND VPWR VPWR _1727_/D sky130_fd_sc_hd__and2_1
X_1655_ _2381_/Q _2378_/Q VGND VGND VPWR VPWR _1655_/X sky130_fd_sc_hd__and2_1
X_1586_ _2445_/Q _1586_/B _2447_/Q _2446_/Q VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__or4b_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _1815_/C _2186_/X _2205_/X _2206_/Y VGND VGND VPWR VPWR _2207_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2138_ _2493_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2138_/X sky130_fd_sc_hd__o31a_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2069_ _2060_/Y _2022_/X _2068_/Y VGND VGND VPWR VPWR _2518_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ _1440_/A VGND VGND VPWR VPWR _2481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1371_ _1371_/A VGND VGND VPWR VPWR _2512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1707_ _1707_/A _1707_/B VGND VGND VPWR VPWR _2394_/D sky130_fd_sc_hd__nor2_1
X_1638_ _2375_/Q _2372_/Q _1637_/B VGND VGND VPWR VPWR _2375_/D sky130_fd_sc_hd__a21o_1
XFILLER_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1569_ _2186_/A VGND VGND VPWR VPWR _1578_/S sky130_fd_sc_hd__clkbuf_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2541_ _2573_/CLK _2541_/D VGND VGND VPWR VPWR _2541_/Q sky130_fd_sc_hd__dfxtp_1
X_2472_ _2503_/CLK _2472_/D _1962_/Y VGND VGND VPWR VPWR _2472_/Q sky130_fd_sc_hd__dfrtp_1
X_1423_ _1423_/A VGND VGND VPWR VPWR _2489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1354_ _2550_/Q _1339_/X _1351_/X _1353_/Y VGND VGND VPWR VPWR _2549_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1285_ _2563_/Q _1261_/X _1282_/X _1284_/Y VGND VGND VPWR VPWR _2562_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1972_ _1974_/A VGND VGND VPWR VPWR _1972_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2524_ _2528_/CLK _2524_/D VGND VGND VPWR VPWR _2524_/Q sky130_fd_sc_hd__dfxtp_1
X_2455_ _2489_/CLK _2455_/D _1941_/Y VGND VGND VPWR VPWR _2455_/Q sky130_fd_sc_hd__dfrtp_1
X_2386_ _2395_/CLK _2386_/D _1855_/Y VGND VGND VPWR VPWR _2386_/Q sky130_fd_sc_hd__dfrtp_1
X_1406_ _2496_/Q _2497_/Q _1406_/S VGND VGND VPWR VPWR _1407_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1337_ _1320_/X _1313_/X _1336_/Y VGND VGND VPWR VPWR _1337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1268_ _1293_/A VGND VGND VPWR VPWR _1268_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1199_ input58/X _1191_/X _1339_/A VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _1243_/Y _2237_/X _2205_/X _2239_/Y VGND VGND VPWR VPWR _2240_/Y sky130_fd_sc_hd__o211ai_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2171_ _2171_/A _2228_/B VGND VGND VPWR VPWR _2171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1955_ _1956_/A VGND VGND VPWR VPWR _1955_/Y sky130_fd_sc_hd__inv_2
X_1886_ _1887_/A VGND VGND VPWR VPWR _1886_/Y sky130_fd_sc_hd__inv_2
X_2507_ _2510_/CLK _2507_/D _2005_/Y VGND VGND VPWR VPWR _2507_/Q sky130_fd_sc_hd__dfrtp_1
X_2438_ _2578_/CLK _2438_/D _1921_/Y VGND VGND VPWR VPWR _2438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2369_ _2601_/CLK _2369_/D _1835_/Y VGND VGND VPWR VPWR _2369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1740_ _1740_/A VGND VGND VPWR VPWR _2404_/D sky130_fd_sc_hd__clkbuf_1
X_1671_ _1631_/X _1673_/C _1673_/D _1673_/B VGND VGND VPWR VPWR _1674_/A sky130_fd_sc_hd__o22a_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2223_ _1254_/Y _2135_/X _2205_/X _2222_/Y VGND VGND VPWR VPWR _2223_/Y sky130_fd_sc_hd__o211ai_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2154_ _1643_/C _2118_/X _2119_/X _2153_/Y VGND VGND VPWR VPWR _2154_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2085_ _1336_/Y _2062_/X _2074_/X _2084_/Y VGND VGND VPWR VPWR _2085_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ _1944_/A VGND VGND VPWR VPWR _1943_/A sky130_fd_sc_hd__buf_2
X_1869_ _1869_/A VGND VGND VPWR VPWR _1869_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1723_ _2410_/Q VGND VGND VPWR VPWR _1727_/C sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2521_/CLK sky130_fd_sc_hd__clkbuf_16
X_1654_ _2379_/Q _2376_/Q _1653_/B VGND VGND VPWR VPWR _2379_/D sky130_fd_sc_hd__a21o_1
X_1585_ _2444_/Q VGND VGND VPWR VPWR _1586_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2229_/A _2469_/Q VGND VGND VPWR VPWR _2206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2137_ _1304_/Y _2135_/X _2119_/X _2136_/Y VGND VGND VPWR VPWR _2137_/Y sky130_fd_sc_hd__o211ai_1
X_2068_ _2061_/Y _2065_/Y _2067_/X VGND VGND VPWR VPWR _2068_/Y sky130_fd_sc_hd__o21ai_2
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1370_ _2512_/Q _2406_/Q _1372_/S VGND VGND VPWR VPWR _1371_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1706_ _1703_/X _1704_/Y _1706_/C _2413_/Q VGND VGND VPWR VPWR _1707_/B sky130_fd_sc_hd__and4bb_1
X_1637_ _1637_/A _1637_/B VGND VGND VPWR VPWR _2374_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1568_ _1568_/A VGND VGND VPWR VPWR _2415_/D sky130_fd_sc_hd__clkbuf_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A VGND VGND VPWR VPWR _2455_/D sky130_fd_sc_hd__clkbuf_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2540_ _2573_/CLK _2540_/D VGND VGND VPWR VPWR _2540_/Q sky130_fd_sc_hd__dfxtp_1
X_2471_ _2504_/CLK _2471_/D _1961_/Y VGND VGND VPWR VPWR _2471_/Q sky130_fd_sc_hd__dfrtp_1
X_1422_ _2489_/Q _2490_/Q _1428_/S VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__mux2_1
X_1353_ _1346_/X _1341_/X _1352_/Y VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1284_ _1268_/X _1263_/X _2171_/A VGND VGND VPWR VPWR _1284_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1971_ _1974_/A VGND VGND VPWR VPWR _1971_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2523_ _2528_/CLK _2523_/D VGND VGND VPWR VPWR _2523_/Q sky130_fd_sc_hd__dfxtp_1
X_2454_ _2489_/CLK _2454_/D _1940_/Y VGND VGND VPWR VPWR _2454_/Q sky130_fd_sc_hd__dfrtp_1
X_1405_ _1405_/A VGND VGND VPWR VPWR _2497_/D sky130_fd_sc_hd__clkbuf_1
X_2385_ _2406_/CLK _2385_/D _1854_/Y VGND VGND VPWR VPWR _2385_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1336_ _2552_/Q VGND VGND VPWR VPWR _1336_/Y sky130_fd_sc_hd__inv_2
Xinput1 wb_rst_i VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1267_ input45/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1198_ _1497_/A VGND VGND VPWR VPWR _1339_/A sky130_fd_sc_hd__buf_4
XFILLER_12_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2170_/A VGND VGND VPWR VPWR _2228_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1954_ _1956_/A VGND VGND VPWR VPWR _1954_/Y sky130_fd_sc_hd__inv_2
X_1885_ _1887_/A VGND VGND VPWR VPWR _1885_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2506_ _2510_/CLK _2506_/D _2004_/Y VGND VGND VPWR VPWR _2506_/Q sky130_fd_sc_hd__dfrtp_1
X_2437_ _2573_/CLK _2437_/D _1918_/Y VGND VGND VPWR VPWR _2437_/Q sky130_fd_sc_hd__dfrtp_4
X_2368_ _2601_/CLK _2368_/D _1834_/Y VGND VGND VPWR VPWR _2368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2299_ input1/X VGND VGND VPWR VPWR _2324_/A sky130_fd_sc_hd__buf_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1319_ _2066_/A VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__clkbuf_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1670_ _2385_/Q _2382_/Q VGND VGND VPWR VPWR _1673_/B sky130_fd_sc_hd__nor2_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2229_/A _2471_/Q VGND VGND VPWR VPWR _2222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2153_ _2187_/A _2463_/Q VGND VGND VPWR VPWR _2153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2084_ _2099_/A _2455_/Q VGND VGND VPWR VPWR _2084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1937_ _1937_/A VGND VGND VPWR VPWR _1937_/Y sky130_fd_sc_hd__inv_2
X_1868_ _1869_/A VGND VGND VPWR VPWR _1868_/Y sky130_fd_sc_hd__inv_2
X_1799_ _2595_/Q _2592_/Q VGND VGND VPWR VPWR _1799_/X sky130_fd_sc_hd__and2_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1722_ _1722_/A VGND VGND VPWR VPWR _1722_/X sky130_fd_sc_hd__clkbuf_4
X_1653_ _1653_/A _1653_/B VGND VGND VPWR VPWR _2378_/D sky130_fd_sc_hd__nor2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1584_/A VGND VGND VPWR VPWR _2408_/D sky130_fd_sc_hd__clkbuf_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2249_/A VGND VGND VPWR VPWR _2205_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2136_ _2144_/A _2461_/Q VGND VGND VPWR VPWR _2136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2067_ _2485_/Q _2066_/X _2016_/X _2056_/X VGND VGND VPWR VPWR _2067_/X sky130_fd_sc_hd__o31a_1
XFILLER_81_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1705_ _1702_/X _2413_/Q _1703_/X _1704_/Y VGND VGND VPWR VPWR _1707_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1636_ _1643_/A _1636_/B _1636_/C _1636_/D VGND VGND VPWR VPWR _1637_/B sky130_fd_sc_hd__nor4_1
X_1567_ input64/X _2415_/Q _1567_/S VGND VGND VPWR VPWR _1568_/A sky130_fd_sc_hd__mux2_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _2455_/Q _2456_/Q _1506_/S VGND VGND VPWR VPWR _1499_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2119_ _2249_/A VGND VGND VPWR VPWR _2119_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2470_ _2503_/CLK _2470_/D _1960_/Y VGND VGND VPWR VPWR _2470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1421_ _1421_/A VGND VGND VPWR VPWR _2490_/D sky130_fd_sc_hd__clkbuf_1
X_1352_ _2549_/Q VGND VGND VPWR VPWR _1352_/Y sky130_fd_sc_hd__inv_2
X_1283_ _2562_/Q VGND VGND VPWR VPWR _2171_/A sky130_fd_sc_hd__inv_2
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2504_/CLK sky130_fd_sc_hd__clkbuf_16
X_1619_ _2371_/Q _2368_/Q VGND VGND VPWR VPWR _1621_/B sky130_fd_sc_hd__nor2_1
X_2599_ _2601_/CLK _2599_/D _2365_/Y VGND VGND VPWR VPWR _2599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1970_ _1974_/A VGND VGND VPWR VPWR _1970_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2522_ _2528_/CLK _2522_/D VGND VGND VPWR VPWR _2522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2453_ _2453_/CLK _2453_/D _1939_/Y VGND VGND VPWR VPWR _2453_/Q sky130_fd_sc_hd__dfrtp_1
X_2384_ _2406_/CLK _2384_/D _1853_/Y VGND VGND VPWR VPWR _2384_/Q sky130_fd_sc_hd__dfrtp_1
X_1404_ _2497_/Q _2498_/Q _1406_/S VGND VGND VPWR VPWR _1405_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1335_ input63/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1335_/X sky130_fd_sc_hd__o21ba_1
Xinput2 wbs_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1266_ _2567_/Q _1261_/X _1262_/X _1265_/Y VGND VGND VPWR VPWR _2566_/D sky130_fd_sc_hd__a22o_1
X_1197_ _2448_/Q VGND VGND VPWR VPWR _1497_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1953_ _1956_/A VGND VGND VPWR VPWR _1953_/Y sky130_fd_sc_hd__inv_2
X_1884_ _1887_/A VGND VGND VPWR VPWR _1884_/Y sky130_fd_sc_hd__inv_2
X_2505_ _2505_/CLK _2505_/D _2003_/Y VGND VGND VPWR VPWR _2505_/Q sky130_fd_sc_hd__dfrtp_1
X_2436_ _2573_/CLK _2436_/D _1917_/Y VGND VGND VPWR VPWR _2436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2367_ _2367_/A VGND VGND VPWR VPWR _2367_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2298_ _2291_/Y _2116_/A _2297_/Y VGND VGND VPWR VPWR _2545_/D sky130_fd_sc_hd__o21ai_1
X_1318_ _1512_/D VGND VGND VPWR VPWR _2066_/A sky130_fd_sc_hd__clkbuf_4
X_1249_ _1242_/X _1237_/X _2228_/A VGND VGND VPWR VPWR _1249_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2264_/A _2236_/B _2430_/Q VGND VGND VPWR VPWR _2221_/Y sky130_fd_sc_hd__nor3b_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2152_ _2238_/A VGND VGND VPWR VPWR _2187_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2083_ _2083_/A _2134_/B _2414_/Q VGND VGND VPWR VPWR _2083_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1936_ _1937_/A VGND VGND VPWR VPWR _1936_/Y sky130_fd_sc_hd__inv_2
X_1867_ _1869_/A VGND VGND VPWR VPWR _1867_/Y sky130_fd_sc_hd__inv_2
Xinput60 wbs_dat_i[3] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1798_ _2593_/Q _2590_/Q _1797_/B VGND VGND VPWR VPWR _2593_/D sky130_fd_sc_hd__a21o_1
X_2419_ _2528_/CLK _2419_/D _1897_/Y VGND VGND VPWR VPWR _2419_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1721_ _2399_/Q _2396_/Q _1720_/B VGND VGND VPWR VPWR _2399_/D sky130_fd_sc_hd__a21o_1
X_1652_ _1648_/X _1649_/Y _1652_/C _2421_/Q VGND VGND VPWR VPWR _1653_/B sky130_fd_sc_hd__and4bb_1
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1583_ input35/X _2408_/Q _1583_/S VGND VGND VPWR VPWR _1584_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2204_/A _2228_/B VGND VGND VPWR VPWR _2204_/Y sky130_fd_sc_hd__nor2_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2135_ _2237_/A VGND VGND VPWR VPWR _2135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2066_ _2066_/A VGND VGND VPWR VPWR _2066_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1919_ _2361_/A VGND VGND VPWR VPWR _1944_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1704_ _2395_/Q _2392_/Q VGND VGND VPWR VPWR _1704_/Y sky130_fd_sc_hd__nor2_1
X_1635_ _1631_/X _1636_/C _1636_/D _1636_/B VGND VGND VPWR VPWR _1637_/A sky130_fd_sc_hd__o22a_1
X_1566_ _1566_/A VGND VGND VPWR VPWR _2416_/D sky130_fd_sc_hd__clkbuf_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1497_/A VGND VGND VPWR VPWR _1506_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2118_ _2186_/A VGND VGND VPWR VPWR _2118_/X sky130_fd_sc_hd__clkbuf_2
X_2049_ _2483_/Q _1346_/A _2016_/X _2246_/A VGND VGND VPWR VPWR _2049_/X sky130_fd_sc_hd__o31a_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1420_ _2490_/Q _2491_/Q _1428_/S VGND VGND VPWR VPWR _1421_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1351_ input60/X _2046_/B _1330_/X VGND VGND VPWR VPWR _1351_/X sky130_fd_sc_hd__o21ba_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1282_ input42/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__o21ba_1
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1618_ _2371_/Q _2368_/Q VGND VGND VPWR VPWR _1621_/D sky130_fd_sc_hd__and2_1
X_2598_ _2601_/CLK _2598_/D _2364_/Y VGND VGND VPWR VPWR _2598_/Q sky130_fd_sc_hd__dfrtp_1
X_1549_ _1549_/A VGND VGND VPWR VPWR _2424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2521_ _2521_/CLK _2521_/D VGND VGND VPWR VPWR _2521_/Q sky130_fd_sc_hd__dfxtp_1
X_2452_ _2453_/CLK _2452_/D _1937_/Y VGND VGND VPWR VPWR _2452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2383_ _2387_/CLK _2383_/D _1852_/Y VGND VGND VPWR VPWR _2383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1403_ _1403_/A VGND VGND VPWR VPWR _2498_/D sky130_fd_sc_hd__clkbuf_1
X_1334_ _2554_/Q _1311_/X _1331_/X _1333_/Y VGND VGND VPWR VPWR _2553_/D sky130_fd_sc_hd__a22o_1
X_1265_ _1242_/X _1263_/X _2204_/A VGND VGND VPWR VPWR _1265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput3 wbs_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1196_ input59/X _1191_/X _1195_/Y VGND VGND VPWR VPWR _2577_/D sky130_fd_sc_hd__o21a_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ _1956_/A VGND VGND VPWR VPWR _1952_/Y sky130_fd_sc_hd__inv_2
X_1883_ _1887_/A VGND VGND VPWR VPWR _1883_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2504_ _2504_/CLK _2504_/D _2002_/Y VGND VGND VPWR VPWR _2504_/Q sky130_fd_sc_hd__dfrtp_1
X_2435_ _2573_/CLK _2435_/D _1916_/Y VGND VGND VPWR VPWR _2435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2366_ _2366_/A VGND VGND VPWR VPWR _2366_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1317_ input66/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1317_/X sky130_fd_sc_hd__o21ba_1
X_2297_ _2292_/Y _2295_/Y _2296_/X VGND VGND VPWR VPWR _2297_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1248_ _2569_/Q VGND VGND VPWR VPWR _2228_/A sky130_fd_sc_hd__inv_2
XFILLER_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1179_ _1179_/A input2/X VGND VGND VPWR VPWR _1182_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2536_/Q VGND VGND VPWR VPWR _2220_/Y sky130_fd_sc_hd__inv_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2151_ _2151_/A _2161_/B VGND VGND VPWR VPWR _2151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2082_ _2520_/Q VGND VGND VPWR VPWR _2082_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1935_ _1937_/A VGND VGND VPWR VPWR _1935_/Y sky130_fd_sc_hd__inv_2
X_1866_ _1869_/A VGND VGND VPWR VPWR _1866_/Y sky130_fd_sc_hd__inv_2
Xinput50 wbs_dat_i[23] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_dat_i[4] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1797_ _1797_/A _1797_/B VGND VGND VPWR VPWR _2592_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2418_ _2555_/CLK _2418_/D _1896_/Y VGND VGND VPWR VPWR _2418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2349_ _2355_/A VGND VGND VPWR VPWR _2354_/A sky130_fd_sc_hd__buf_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1720_ _1720_/A _1720_/B VGND VGND VPWR VPWR _2398_/D sky130_fd_sc_hd__nor2_1
X_1651_ _2546_/Q VGND VGND VPWR VPWR _1652_/C sky130_fd_sc_hd__clkbuf_2
X_1582_ _1582_/A VGND VGND VPWR VPWR _2409_/D sky130_fd_sc_hd__clkbuf_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2246_/A VGND VGND VPWR VPWR _2203_/X sky130_fd_sc_hd__clkbuf_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _2194_/A _2134_/B _2420_/Q VGND VGND VPWR VPWR _2134_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2065_ _1347_/Y _2062_/X _2030_/X _2064_/Y VGND VGND VPWR VPWR _2065_/Y sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2446_/CLK sky130_fd_sc_hd__clkbuf_16
X_1918_ _1918_/A VGND VGND VPWR VPWR _1918_/Y sky130_fd_sc_hd__inv_2
X_1849_ _1850_/A VGND VGND VPWR VPWR _1849_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1703_ _2395_/Q _2392_/Q VGND VGND VPWR VPWR _1703_/X sky130_fd_sc_hd__and2_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1634_ _2375_/Q _2372_/Q VGND VGND VPWR VPWR _1636_/B sky130_fd_sc_hd__nor2_1
X_1565_ input65/X _2416_/Q _1567_/S VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__mux2_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1496_/A VGND VGND VPWR VPWR _2456_/D sky130_fd_sc_hd__clkbuf_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2117_ _2117_/A _2161_/B VGND VGND VPWR VPWR _2117_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2048_ _1727_/C _1583_/S _2030_/X _2047_/Y VGND VGND VPWR VPWR _2048_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_54_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1350_ _2170_/A VGND VGND VPWR VPWR _2046_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ _2564_/Q _1261_/X _1278_/X _1280_/Y VGND VGND VPWR VPWR _2563_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1617_ _2425_/Q VGND VGND VPWR VPWR _1621_/C sky130_fd_sc_hd__clkinv_2
X_2597_ _2597_/CLK _2597_/D _2363_/Y VGND VGND VPWR VPWR _2597_/Q sky130_fd_sc_hd__dfrtp_1
X_1548_ input42/X _2424_/Q _1556_/S VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1479_ _1479_/A VGND VGND VPWR VPWR _2464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2536_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2520_ _2520_/CLK _2520_/D VGND VGND VPWR VPWR _2520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2451_ _2484_/CLK _2451_/D _1936_/Y VGND VGND VPWR VPWR _2451_/Q sky130_fd_sc_hd__dfrtp_1
X_1402_ _2498_/Q _2499_/Q _1406_/S VGND VGND VPWR VPWR _1403_/A sky130_fd_sc_hd__mux2_1
X_2382_ _2406_/CLK _2382_/D _1850_/Y VGND VGND VPWR VPWR _2382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1333_ _1320_/X _1313_/X _2091_/A VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1264_ _2566_/Q VGND VGND VPWR VPWR _2204_/A sky130_fd_sc_hd__inv_2
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 wbs_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_1195_ _2292_/A _1191_/X _1194_/X VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1951_ _1975_/A VGND VGND VPWR VPWR _1956_/A sky130_fd_sc_hd__buf_2
X_1882_ _1882_/A VGND VGND VPWR VPWR _1887_/A sky130_fd_sc_hd__buf_4
X_2503_ _2503_/CLK _2503_/D _2001_/Y VGND VGND VPWR VPWR _2503_/Q sky130_fd_sc_hd__dfrtp_1
X_2434_ _2539_/CLK _2434_/D _1915_/Y VGND VGND VPWR VPWR _2434_/Q sky130_fd_sc_hd__dfrtp_1
X_2365_ _2366_/A VGND VGND VPWR VPWR _2365_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1316_ _2557_/Q _1311_/X _1312_/X _1315_/Y VGND VGND VPWR VPWR _2556_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2296_ _2512_/Q _2066_/A _2165_/A _2032_/X VGND VGND VPWR VPWR _2296_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1247_ input50/X _1246_/X _1224_/X VGND VGND VPWR VPWR _1247_/X sky130_fd_sc_hd__o21ba_1
X_1178_ _1178_/A _1178_/B VGND VGND VPWR VPWR _2028_/B sky130_fd_sc_hd__nor2_8
XFILLER_64_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2150_ _2528_/Q VGND VGND VPWR VPWR _2150_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2081_ _2070_/Y _2071_/X _2080_/Y VGND VGND VPWR VPWR _2519_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1934_ _1937_/A VGND VGND VPWR VPWR _1934_/Y sky130_fd_sc_hd__inv_2
X_1865_ _1869_/A VGND VGND VPWR VPWR _1865_/Y sky130_fd_sc_hd__inv_2
Xinput40 wbs_dat_i[14] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 wbs_dat_i[24] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_dat_i[5] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
X_1796_ _1828_/A _1796_/B _1796_/C _1796_/D VGND VGND VPWR VPWR _1797_/B sky130_fd_sc_hd__nor4_1
X_2417_ _2521_/CLK _2417_/D _1894_/Y VGND VGND VPWR VPWR _2417_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2348_ _2348_/A VGND VGND VPWR VPWR _2348_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2279_ _2294_/A _2478_/Q VGND VGND VPWR VPWR _2279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1650_ _1647_/X _2421_/Q _1648_/X _1649_/Y VGND VGND VPWR VPWR _1653_/A sky130_fd_sc_hd__o2bb2a_1
X_1581_ input46/X _2409_/Q _1583_/S VGND VGND VPWR VPWR _1582_/A sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2534_/Q VGND VGND VPWR VPWR _2202_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _2526_/Q VGND VGND VPWR VPWR _2133_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2064_ _2099_/A _2453_/Q VGND VGND VPWR VPWR _2064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1917_ _1918_/A VGND VGND VPWR VPWR _1917_/Y sky130_fd_sc_hd__inv_2
X_1848_ _1850_/A VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__inv_2
X_1779_ _2587_/Q _2584_/Q _1778_/B VGND VGND VPWR VPWR _2587_/D sky130_fd_sc_hd__a21o_1
XFILLER_1_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1702_ _1747_/A VGND VGND VPWR VPWR _1702_/X sky130_fd_sc_hd__buf_2
XFILLER_8_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1633_ _2375_/Q _2372_/Q VGND VGND VPWR VPWR _1636_/D sky130_fd_sc_hd__and2_1
X_1564_ _1564_/A VGND VGND VPWR VPWR _2417_/D sky130_fd_sc_hd__clkbuf_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _2456_/Q _2457_/Q _1495_/S VGND VGND VPWR VPWR _1496_/A sky130_fd_sc_hd__mux2_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2116_ _2116_/A VGND VGND VPWR VPWR _2116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2047_ _2054_/A _2451_/Q VGND VGND VPWR VPWR _2047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2453_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _1268_/X _1263_/X _2178_/A VGND VGND VPWR VPWR _1280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2596_ _2601_/CLK _2596_/D _2362_/Y VGND VGND VPWR VPWR _2596_/Q sky130_fd_sc_hd__dfrtp_1
X_1616_ _1672_/A VGND VGND VPWR VPWR _1828_/A sky130_fd_sc_hd__buf_2
X_1547_ _1558_/A VGND VGND VPWR VPWR _1556_/S sky130_fd_sc_hd__buf_2
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1478_ _2464_/Q _2465_/Q _1484_/S VGND VGND VPWR VPWR _1479_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2450_ _2484_/CLK _2450_/D _1935_/Y VGND VGND VPWR VPWR _2450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1401_ _1401_/A VGND VGND VPWR VPWR _2499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2381_ _2387_/CLK _2381_/D _1849_/Y VGND VGND VPWR VPWR _2381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1332_ _2553_/Q VGND VGND VPWR VPWR _2091_/A sky130_fd_sc_hd__inv_2
XFILLER_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1263_ _2024_/B VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 wbs_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_1194_ _1589_/A VGND VGND VPWR VPWR _1194_/X sky130_fd_sc_hd__buf_8
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2579_ _2587_/CLK _2579_/D _2341_/Y VGND VGND VPWR VPWR _2579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ input1/X VGND VGND VPWR VPWR _1975_/A sky130_fd_sc_hd__buf_2
X_1881_ _1881_/A VGND VGND VPWR VPWR _1881_/Y sky130_fd_sc_hd__inv_2
X_2502_ _2503_/CLK _2502_/D _1999_/Y VGND VGND VPWR VPWR _2502_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2433_ _2539_/CLK _2433_/D _1914_/Y VGND VGND VPWR VPWR _2433_/Q sky130_fd_sc_hd__dfrtp_4
X_2364_ _2366_/A VGND VGND VPWR VPWR _2364_/Y sky130_fd_sc_hd__inv_2
X_1315_ _1293_/X _1313_/X _2117_/A VGND VGND VPWR VPWR _1315_/Y sky130_fd_sc_hd__o21ai_1
X_2295_ _2293_/Y _2186_/X _2074_/A _2294_/Y VGND VGND VPWR VPWR _2295_/Y sky130_fd_sc_hd__o211ai_2
X_1246_ _1297_/A VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1177_ _1177_/A _1177_/B _1177_/C _1177_/D VGND VGND VPWR VPWR _1178_/B sky130_fd_sc_hd__nand4_4
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2080_ _2073_/Y _2076_/Y _2079_/X VGND VGND VPWR VPWR _2080_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1933_ _1937_/A VGND VGND VPWR VPWR _1933_/Y sky130_fd_sc_hd__inv_2
Xinput30 wbs_adr_i[6] VGND VGND VPWR VPWR _1166_/B sky130_fd_sc_hd__clkbuf_1
X_1864_ _1882_/A VGND VGND VPWR VPWR _1869_/A sky130_fd_sc_hd__buf_2
Xinput63 wbs_dat_i[6] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_dat_i[15] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 wbs_dat_i[25] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
X_1795_ _1722_/X _1796_/C _1796_/D _1796_/B VGND VGND VPWR VPWR _1797_/A sky130_fd_sc_hd__o22a_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2416_ _2555_/CLK _2416_/D _1893_/Y VGND VGND VPWR VPWR _2416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2347_ _2348_/A VGND VGND VPWR VPWR _2347_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2278_ _2285_/A _2285_/B _2437_/Q VGND VGND VPWR VPWR _2278_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ input53/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1229_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1580_ _2186_/A VGND VGND VPWR VPWR _1583_/S sky130_fd_sc_hd__clkbuf_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2193_/Y _2160_/X _2200_/Y VGND VGND VPWR VPWR _2533_/D sky130_fd_sc_hd__o21ai_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2132_ _2126_/Y _2116_/X _2131_/Y VGND VGND VPWR VPWR _2525_/D sky130_fd_sc_hd__o21ai_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2063_ _2247_/A VGND VGND VPWR VPWR _2099_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1916_ _1918_/A VGND VGND VPWR VPWR _1916_/Y sky130_fd_sc_hd__inv_2
X_1847_ _1850_/A VGND VGND VPWR VPWR _1847_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2510_/CLK sky130_fd_sc_hd__clkbuf_16
X_1778_ _1778_/A _1778_/B VGND VGND VPWR VPWR _2586_/D sky130_fd_sc_hd__nor2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1701_ _2393_/Q _2390_/Q _1700_/B VGND VGND VPWR VPWR _2393_/D sky130_fd_sc_hd__a21o_1
X_1632_ _2423_/Q VGND VGND VPWR VPWR _1636_/C sky130_fd_sc_hd__clkinv_2
X_1563_ input66/X _2417_/Q _1567_/S VGND VGND VPWR VPWR _1564_/A sky130_fd_sc_hd__mux2_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1494_/A VGND VGND VPWR VPWR _2457_/D sky130_fd_sc_hd__clkbuf_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2115_ _2524_/Q VGND VGND VPWR VPWR _2115_/Y sky130_fd_sc_hd__inv_2
X_2046_ _2046_/A _2046_/B VGND VGND VPWR VPWR _2046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1615_ _1615_/A VGND VGND VPWR VPWR _2447_/D sky130_fd_sc_hd__clkbuf_1
X_2595_ _2597_/CLK _2595_/D _2360_/Y VGND VGND VPWR VPWR _2595_/Q sky130_fd_sc_hd__dfrtp_1
X_1546_ _1546_/A VGND VGND VPWR VPWR _2425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1477_ _1477_/A VGND VGND VPWR VPWR _2465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2029_ _2249_/A VGND VGND VPWR VPWR _2074_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ _2499_/Q _2500_/Q _1406_/S VGND VGND VPWR VPWR _1401_/A sky130_fd_sc_hd__mux2_1
X_2380_ _2387_/CLK _2380_/D _1848_/Y VGND VGND VPWR VPWR _2380_/Q sky130_fd_sc_hd__dfrtp_1
X_1331_ input64/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__o21ba_1
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1262_ input47/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__o21ba_1
Xinput6 wbs_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
X_1193_ _2448_/Q VGND VGND VPWR VPWR _1589_/A sky130_fd_sc_hd__buf_6
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2578_ _2578_/CLK _2578_/D _2340_/Y VGND VGND VPWR VPWR _2578_/Q sky130_fd_sc_hd__dfrtp_1
X_1529_ _1529_/A VGND VGND VPWR VPWR _2433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1880_ _1881_/A VGND VGND VPWR VPWR _1880_/Y sky130_fd_sc_hd__inv_2
X_2501_ _2505_/CLK _2501_/D _1998_/Y VGND VGND VPWR VPWR _2501_/Q sky130_fd_sc_hd__dfrtp_1
X_2432_ _2539_/CLK _2432_/D _1912_/Y VGND VGND VPWR VPWR _2432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2363_ _2366_/A VGND VGND VPWR VPWR _2363_/Y sky130_fd_sc_hd__inv_2
X_1314_ _2556_/Q VGND VGND VPWR VPWR _2117_/A sky130_fd_sc_hd__inv_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2294_ _2294_/A _2480_/Q VGND VGND VPWR VPWR _2294_/Y sky130_fd_sc_hd__nand2_1
X_1245_ _2571_/Q _1233_/X _1241_/X _1244_/Y VGND VGND VPWR VPWR _2570_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1176_ _1176_/A _1176_/B VGND VGND VPWR VPWR _1177_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1932_ _1944_/A VGND VGND VPWR VPWR _1937_/A sky130_fd_sc_hd__buf_2
X_1863_ _1863_/A VGND VGND VPWR VPWR _1863_/Y sky130_fd_sc_hd__inv_2
Xinput31 wbs_adr_i[7] VGND VGND VPWR VPWR _1166_/A sky130_fd_sc_hd__clkbuf_1
Xinput20 wbs_adr_i[26] VGND VGND VPWR VPWR _1176_/B sky130_fd_sc_hd__clkbuf_1
Xinput53 wbs_dat_i[26] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_dat_i[7] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
Xinput42 wbs_dat_i[16] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
X_1794_ _2593_/Q _2590_/Q VGND VGND VPWR VPWR _1796_/B sky130_fd_sc_hd__nor2_1
X_2415_ _2521_/CLK _2415_/D _1892_/Y VGND VGND VPWR VPWR _2415_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2346_ _2348_/A VGND VGND VPWR VPWR _2346_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2277_ _2543_/Q VGND VGND VPWR VPWR _2277_/Y sky130_fd_sc_hd__inv_2
X_1228_ _2574_/Q _1209_/X _1225_/X _1227_/Y VGND VGND VPWR VPWR _2573_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2194_/Y _2197_/Y _2199_/X VGND VGND VPWR VPWR _2200_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2131_ _2127_/Y _2129_/Y _2130_/X VGND VGND VPWR VPWR _2131_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2062_ _2170_/A VGND VGND VPWR VPWR _2062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1915_ _1918_/A VGND VGND VPWR VPWR _1915_/Y sky130_fd_sc_hd__inv_2
X_1846_ _1850_/A VGND VGND VPWR VPWR _1846_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1777_ _1777_/A _1777_/B _1777_/C _1777_/D VGND VGND VPWR VPWR _1778_/B sky130_fd_sc_hd__nor4_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2329_/A VGND VGND VPWR VPWR _2329_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1700_ _1700_/A _1700_/B VGND VGND VPWR VPWR _2392_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1631_ _1672_/A VGND VGND VPWR VPWR _1631_/X sky130_fd_sc_hd__buf_2
X_1562_ _1562_/A VGND VGND VPWR VPWR _2418_/D sky130_fd_sc_hd__clkbuf_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _2457_/Q _2458_/Q _1495_/S VGND VGND VPWR VPWR _1494_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2114_ _2105_/Y _2071_/X _2113_/Y VGND VGND VPWR VPWR _2523_/D sky130_fd_sc_hd__o21ai_1
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2045_ _2516_/Q VGND VGND VPWR VPWR _2045_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1829_ _1829_/A _1829_/B VGND VGND VPWR VPWR _2368_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1614_ _1614_/A _1614_/B _1614_/C VGND VGND VPWR VPWR _1615_/A sky130_fd_sc_hd__and3_1
X_2594_ _2597_/CLK _2594_/D _2359_/Y VGND VGND VPWR VPWR _2594_/Q sky130_fd_sc_hd__dfrtp_1
X_1545_ input43/X _2425_/Q _1545_/S VGND VGND VPWR VPWR _1546_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1476_ _2465_/Q _2466_/Q _1484_/S VGND VGND VPWR VPWR _1477_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2028_ _2213_/A _2028_/B _2028_/C _2028_/D VGND VGND VPWR VPWR _2249_/A sky130_fd_sc_hd__nand4_4
XFILLER_23_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1330_ _1374_/A VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1261_ _1608_/B VGND VGND VPWR VPWR _1261_/X sky130_fd_sc_hd__clkbuf_2
Xinput7 wbs_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
X_1192_ _2577_/Q VGND VGND VPWR VPWR _2292_/A sky130_fd_sc_hd__inv_2
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2577_ _2577_/CLK _2577_/D _2339_/Y VGND VGND VPWR VPWR _2577_/Q sky130_fd_sc_hd__dfrtp_1
X_1528_ input52/X _2433_/Q _1534_/S VGND VGND VPWR VPWR _1529_/A sky130_fd_sc_hd__mux2_1
X_1459_ _1459_/A VGND VGND VPWR VPWR _2473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2500_ _2503_/CLK _2500_/D _1997_/Y VGND VGND VPWR VPWR _2500_/Q sky130_fd_sc_hd__dfrtp_1
X_2431_ _2568_/CLK _2431_/D _1911_/Y VGND VGND VPWR VPWR _2431_/Q sky130_fd_sc_hd__dfrtp_1
X_2362_ _2366_/A VGND VGND VPWR VPWR _2362_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1313_ _2024_/B VGND VGND VPWR VPWR _1313_/X sky130_fd_sc_hd__clkbuf_2
X_2293_ _2439_/Q VGND VGND VPWR VPWR _2293_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1244_ _1242_/X _1237_/X _1243_/Y VGND VGND VPWR VPWR _1244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1175_ _1175_/A _1175_/B VGND VGND VPWR VPWR _1177_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2589_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1931_ _1931_/A VGND VGND VPWR VPWR _1931_/Y sky130_fd_sc_hd__inv_2
X_1862_ _1863_/A VGND VGND VPWR VPWR _1862_/Y sky130_fd_sc_hd__inv_2
Xinput10 wbs_adr_i[17] VGND VGND VPWR VPWR _1183_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[27] VGND VGND VPWR VPWR _1176_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 wbs_dat_i[27] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
Xinput32 wbs_adr_i[8] VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_dat_i[17] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
X_1793_ _2593_/Q _2590_/Q VGND VGND VPWR VPWR _1796_/D sky130_fd_sc_hd__and2_1
Xinput65 wbs_dat_i[8] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_1
X_2414_ _2520_/CLK _2414_/D _1891_/Y VGND VGND VPWR VPWR _2414_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2345_ _2348_/A VGND VGND VPWR VPWR _2345_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2276_ _2270_/Y _2246_/X _2275_/Y VGND VGND VPWR VPWR _2542_/D sky130_fd_sc_hd__o21ai_1
XFILLER_84_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1227_ _1212_/X _1214_/X _1226_/Y VGND VGND VPWR VPWR _1227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ _2492_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2130_/X sky130_fd_sc_hd__o31a_1
X_2061_ _2083_/A _2061_/B _2412_/Q VGND VGND VPWR VPWR _2061_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1914_ _1918_/A VGND VGND VPWR VPWR _1914_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1845_ _2367_/A VGND VGND VPWR VPWR _1850_/A sky130_fd_sc_hd__buf_2
X_1776_ _1722_/X _1777_/C _1777_/D _1777_/B VGND VGND VPWR VPWR _1778_/A sky130_fd_sc_hd__o22a_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2328_ _2329_/A VGND VGND VPWR VPWR _2328_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2259_ _1777_/C _2186_/X _2249_/X _2258_/Y VGND VGND VPWR VPWR _2259_/Y sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2496_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ _2373_/Q _2370_/Q _1629_/B VGND VGND VPWR VPWR _2373_/D sky130_fd_sc_hd__a21o_1
X_1561_ input36/X _2418_/Q _1567_/S VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__mux2_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1492_/A VGND VGND VPWR VPWR _2458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2113_ _2107_/Y _2110_/Y _2112_/X VGND VGND VPWR VPWR _2113_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2044_ _2036_/Y _2022_/X _2043_/Y VGND VGND VPWR VPWR _2515_/D sky130_fd_sc_hd__o21ai_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1828_ _1828_/A _1828_/B _1828_/C _1828_/D VGND VGND VPWR VPWR _1829_/B sky130_fd_sc_hd__nor4_1
X_1759_ _1759_/A _1759_/B VGND VGND VPWR VPWR _2580_/D sky130_fd_sc_hd__nor2_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1613_ _2445_/Q _1586_/B _2446_/Q _1606_/C _2447_/Q VGND VGND VPWR VPWR _1614_/B
+ sky130_fd_sc_hd__a41o_1
X_2593_ _2593_/CLK _2593_/D _2358_/Y VGND VGND VPWR VPWR _2593_/Q sky130_fd_sc_hd__dfrtp_1
X_1544_ _1544_/A VGND VGND VPWR VPWR _2426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1475_ _1486_/A VGND VGND VPWR VPWR _1484_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2027_ _2294_/A _2449_/Q VGND VGND VPWR VPWR _2027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1260_ _2568_/Q _1233_/X _1257_/X _1259_/Y VGND VGND VPWR VPWR _2567_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 wbs_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
X_1191_ _2237_/A VGND VGND VPWR VPWR _1191_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2576_ _2577_/CLK _2576_/D _2338_/Y VGND VGND VPWR VPWR _2576_/Q sky130_fd_sc_hd__dfrtp_1
X_1527_ _1527_/A VGND VGND VPWR VPWR _2434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1458_ _2473_/Q _2474_/Q _1462_/S VGND VGND VPWR VPWR _1459_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1389_ _2504_/Q _2505_/Q _1395_/S VGND VGND VPWR VPWR _1390_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2430_ _2568_/CLK _2430_/D _1910_/Y VGND VGND VPWR VPWR _2430_/Q sky130_fd_sc_hd__dfrtp_4
X_2361_ _2361_/A VGND VGND VPWR VPWR _2366_/A sky130_fd_sc_hd__buf_2
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1312_ input36/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1312_/X sky130_fd_sc_hd__o21ba_1
X_2292_ _2292_/A _2292_/B VGND VGND VPWR VPWR _2292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ _2570_/Q VGND VGND VPWR VPWR _1243_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1174_ _1174_/A _1174_/B VGND VGND VPWR VPWR _1177_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2559_ _2560_/CLK _2559_/D _2316_/Y VGND VGND VPWR VPWR _2559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ _1931_/A VGND VGND VPWR VPWR _1930_/Y sky130_fd_sc_hd__inv_2
X_1861_ _1863_/A VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__inv_2
Xinput11 wbs_adr_i[18] VGND VGND VPWR VPWR _1184_/B sky130_fd_sc_hd__clkbuf_1
Xinput22 wbs_adr_i[28] VGND VGND VPWR VPWR _1172_/B sky130_fd_sc_hd__clkbuf_1
X_1792_ _2431_/Q VGND VGND VPWR VPWR _1796_/C sky130_fd_sc_hd__clkinv_2
Xinput55 wbs_dat_i[28] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_1
Xinput33 wbs_adr_i[9] VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_dat_i[18] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput66 wbs_dat_i[9] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2413_ _2520_/CLK _2413_/D _1890_/Y VGND VGND VPWR VPWR _2413_/Q sky130_fd_sc_hd__dfrtp_4
X_2344_ _2348_/A VGND VGND VPWR VPWR _2344_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ _2271_/Y _2273_/Y _2274_/X VGND VGND VPWR VPWR _2275_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1226_ _2573_/Q VGND VGND VPWR VPWR _1226_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2060_ _2518_/Q VGND VGND VPWR VPWR _2060_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1913_ _1913_/A VGND VGND VPWR VPWR _1918_/A sky130_fd_sc_hd__buf_2
X_1844_ _1844_/A VGND VGND VPWR VPWR _1844_/Y sky130_fd_sc_hd__inv_2
X_1775_ _2587_/Q _2584_/Q VGND VGND VPWR VPWR _1777_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2327_ _2329_/A VGND VGND VPWR VPWR _2327_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2258_ _2272_/A _2475_/Q VGND VGND VPWR VPWR _2258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1209_ _1608_/B VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2189_ _2231_/A VGND VGND VPWR VPWR _2189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1560_ _1560_/A VGND VGND VPWR VPWR _2419_/D sky130_fd_sc_hd__clkbuf_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _2458_/Q _2459_/Q _1495_/S VGND VGND VPWR VPWR _1492_/A sky130_fd_sc_hd__mux2_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2112_ _2490_/Q _2111_/X _2078_/X _2101_/X VGND VGND VPWR VPWR _2112_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2043_ _2038_/Y _2040_/Y _2042_/X VGND VGND VPWR VPWR _2043_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1827_ _1722_/X _1828_/C _1828_/D _1828_/B VGND VGND VPWR VPWR _1829_/A sky130_fd_sc_hd__o22a_1
X_1758_ _1754_/X _1755_/Y _1789_/C _2437_/Q VGND VGND VPWR VPWR _1759_/B sky130_fd_sc_hd__and4bb_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1689_ _2415_/Q VGND VGND VPWR VPWR _1693_/C sky130_fd_sc_hd__inv_2
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1612_ _2447_/Q _2446_/Q _1612_/C VGND VGND VPWR VPWR _1614_/A sky130_fd_sc_hd__nand3_1
X_2592_ _2593_/CLK _2592_/D _2357_/Y VGND VGND VPWR VPWR _2592_/Q sky130_fd_sc_hd__dfrtp_1
X_1543_ input44/X _2426_/Q _1545_/S VGND VGND VPWR VPWR _1544_/A sky130_fd_sc_hd__mux2_1
X_1474_ _1474_/A VGND VGND VPWR VPWR _2466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2026_ _2026_/A VGND VGND VPWR VPWR _2294_/A sky130_fd_sc_hd__buf_2
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1190_ _1324_/A VGND VGND VPWR VPWR _2237_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput9 wbs_adr_i[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2575_ _2575_/CLK _2575_/D _2336_/Y VGND VGND VPWR VPWR _2575_/Q sky130_fd_sc_hd__dfrtp_1
X_1526_ input53/X _2434_/Q _1534_/S VGND VGND VPWR VPWR _1527_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1457_ _1457_/A VGND VGND VPWR VPWR _2474_/D sky130_fd_sc_hd__clkbuf_1
X_1388_ _1388_/A VGND VGND VPWR VPWR _2505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2009_ _2011_/A VGND VGND VPWR VPWR _2009_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2360_ _2360_/A VGND VGND VPWR VPWR _2360_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2291_ _2545_/Q VGND VGND VPWR VPWR _2291_/Y sky130_fd_sc_hd__inv_2
X_1311_ _1339_/A VGND VGND VPWR VPWR _1311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1242_ _1293_/A VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1173_ _1173_/A _1173_/B VGND VGND VPWR VPWR _1177_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2573_/CLK sky130_fd_sc_hd__clkbuf_16
X_2558_ _2560_/CLK _2558_/D _2315_/Y VGND VGND VPWR VPWR _2558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2489_ _2489_/CLK _2489_/D _1984_/Y VGND VGND VPWR VPWR _2489_/Q sky130_fd_sc_hd__dfrtp_1
X_1509_ _1509_/A VGND VGND VPWR VPWR _2450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _1863_/A VGND VGND VPWR VPWR _1860_/Y sky130_fd_sc_hd__inv_2
X_1791_ _2591_/Q _2588_/Q _1790_/B VGND VGND VPWR VPWR _2591_/D sky130_fd_sc_hd__a21o_1
Xinput12 wbs_adr_i[19] VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 wbs_dat_i[19] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 wbs_cyc_i VGND VGND VPWR VPWR _1165_/B sky130_fd_sc_hd__clkbuf_1
Xinput23 wbs_adr_i[29] VGND VGND VPWR VPWR _1172_/A sky130_fd_sc_hd__clkbuf_1
Xinput67 wbs_stb_i VGND VGND VPWR VPWR _1165_/A sky130_fd_sc_hd__clkbuf_1
Xinput56 wbs_dat_i[29] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2412_ _2549_/CLK _2412_/D _1887_/Y VGND VGND VPWR VPWR _2412_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2343_ _2355_/A VGND VGND VPWR VPWR _2348_/A sky130_fd_sc_hd__buf_2
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2274_ _2509_/Q _2241_/X _2252_/X _2032_/X VGND VGND VPWR VPWR _2274_/X sky130_fd_sc_hd__o31a_1
X_1225_ input54/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__o21ba_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1989_ _1993_/A VGND VGND VPWR VPWR _1989_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _1912_/A VGND VGND VPWR VPWR _1912_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1843_ _1844_/A VGND VGND VPWR VPWR _1843_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1774_ _2587_/Q _2584_/Q VGND VGND VPWR VPWR _1777_/D sky130_fd_sc_hd__and2_1
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2329_/A VGND VGND VPWR VPWR _2326_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _2257_/A _2292_/B VGND VGND VPWR VPWR _2257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1208_ _1497_/A VGND VGND VPWR VPWR _1608_/B sky130_fd_sc_hd__buf_4
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2188_ _1828_/C _2186_/X _2162_/X _2187_/Y VGND VGND VPWR VPWR _2188_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1490_/A VGND VGND VPWR VPWR _2459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2111_ _2241_/A VGND VGND VPWR VPWR _2111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2042_ _2482_/Q _1346_/A _2016_/X _2246_/A VGND VGND VPWR VPWR _2042_/X sky130_fd_sc_hd__o31a_1
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1826_ _2369_/Q _2600_/Q VGND VGND VPWR VPWR _1828_/B sky130_fd_sc_hd__nor2_1
X_1757_ _2546_/Q VGND VGND VPWR VPWR _1789_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1688_ _2389_/Q _2386_/Q _1687_/B VGND VGND VPWR VPWR _2389_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2311_/A VGND VGND VPWR VPWR _2309_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1611_ _2446_/Q _1612_/C _1610_/Y VGND VGND VPWR VPWR _2446_/D sky130_fd_sc_hd__a21oi_1
X_2591_ _2593_/CLK _2591_/D _2356_/Y VGND VGND VPWR VPWR _2591_/Q sky130_fd_sc_hd__dfrtp_1
X_1542_ _1542_/A VGND VGND VPWR VPWR _2427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1473_ _2466_/Q _2467_/Q _1473_/S VGND VGND VPWR VPWR _1474_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ _2237_/A VGND VGND VPWR VPWR _2292_/B sky130_fd_sc_hd__buf_4
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1809_ _1809_/A _1809_/B VGND VGND VPWR VPWR _2596_/D sky130_fd_sc_hd__nor2_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2574_ _2575_/CLK _2574_/D _2335_/Y VGND VGND VPWR VPWR _2574_/Q sky130_fd_sc_hd__dfrtp_1
X_1525_ _1558_/A VGND VGND VPWR VPWR _1534_/S sky130_fd_sc_hd__buf_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1456_ _2474_/Q _2475_/Q _1462_/S VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1387_ _2505_/Q _2506_/Q _1395_/S VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2008_ _2011_/A VGND VGND VPWR VPWR _2008_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2290_ _2284_/Y _2116_/A _2289_/Y VGND VGND VPWR VPWR _2544_/D sky130_fd_sc_hd__o21ai_1
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1310_ _2558_/Q _1286_/X _1307_/X _1309_/Y VGND VGND VPWR VPWR _2557_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1241_ input51/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__o21ba_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1172_ _1172_/A _1172_/B _1172_/C VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__nand3_2
XFILLER_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 _2522_/Q VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_2557_ _2560_/CLK _2557_/D _2314_/Y VGND VGND VPWR VPWR _2557_/Q sky130_fd_sc_hd__dfrtp_1
X_2488_ _2495_/CLK _2488_/D _1983_/Y VGND VGND VPWR VPWR _2488_/Q sky130_fd_sc_hd__dfrtp_1
X_1508_ _2450_/Q _2451_/Q _1589_/A VGND VGND VPWR VPWR _1509_/A sky130_fd_sc_hd__mux2_1
X_1439_ _2481_/Q _2482_/Q _1439_/S VGND VGND VPWR VPWR _1440_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1790_ _1790_/A _1790_/B VGND VGND VPWR VPWR _2590_/D sky130_fd_sc_hd__nor2_1
Xinput13 wbs_adr_i[1] VGND VGND VPWR VPWR _1179_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 wbs_adr_i[2] VGND VGND VPWR VPWR _1200_/A sky130_fd_sc_hd__buf_2
Xinput46 wbs_dat_i[1] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 wbs_dat_i[0] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_2
Xinput57 wbs_dat_i[2] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput68 wbs_we_i VGND VGND VPWR VPWR _2012_/B sky130_fd_sc_hd__clkbuf_1
X_2411_ _2549_/CLK _2411_/D _1886_/Y VGND VGND VPWR VPWR _2411_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2342_ _2342_/A VGND VGND VPWR VPWR _2342_/Y sky130_fd_sc_hd__inv_2
X_2273_ _1221_/Y _2237_/X _2249_/X _2272_/Y VGND VGND VPWR VPWR _2273_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ _1589_/A VGND VGND VPWR VPWR _1224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1988_ _2006_/A VGND VGND VPWR VPWR _1993_/A sky130_fd_sc_hd__buf_2
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ _1912_/A VGND VGND VPWR VPWR _1911_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1842_ _1844_/A VGND VGND VPWR VPWR _1842_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1773_ _2434_/Q VGND VGND VPWR VPWR _1777_/C sky130_fd_sc_hd__inv_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2329_/A VGND VGND VPWR VPWR _2325_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _2540_/Q VGND VGND VPWR VPWR _2256_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1207_ _1293_/A _2061_/B _1206_/Y VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2187_ _2187_/A _2467_/Q VGND VGND VPWR VPWR _2187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2406_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2110_ _1321_/Y _2062_/X _2074_/X _2109_/Y VGND VGND VPWR VPWR _2110_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2041_ _2146_/A VGND VGND VPWR VPWR _2246_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1825_ _2369_/Q _2600_/Q VGND VGND VPWR VPWR _1828_/D sky130_fd_sc_hd__and2_1
X_1756_ _1747_/X _2437_/Q _1754_/X _1755_/Y VGND VGND VPWR VPWR _1759_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1687_ _1687_/A _1687_/B VGND VGND VPWR VPWR _2388_/D sky130_fd_sc_hd__nor2_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2311_/A VGND VGND VPWR VPWR _2308_/Y sky130_fd_sc_hd__inv_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ _2272_/A _2473_/Q VGND VGND VPWR VPWR _2239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1610_ _2446_/Q _1612_/C _1588_/X _1586_/X _1614_/C VGND VGND VPWR VPWR _1610_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2590_ _2593_/CLK _2590_/D _2354_/Y VGND VGND VPWR VPWR _2590_/Q sky130_fd_sc_hd__dfrtp_1
X_1541_ input45/X _2427_/Q _1545_/S VGND VGND VPWR VPWR _1542_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1472_ _1472_/A VGND VGND VPWR VPWR _2467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2024_ _2285_/A _2024_/B _2408_/Q VGND VGND VPWR VPWR _2024_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1808_ _1805_/X _1806_/Y _1821_/C _2429_/Q VGND VGND VPWR VPWR _1809_/B sky130_fd_sc_hd__and4bb_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1739_ _1737_/X _2405_/D VGND VGND VPWR VPWR _1740_/A sky130_fd_sc_hd__and2b_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2573_ _2573_/CLK _2573_/D _2334_/Y VGND VGND VPWR VPWR _2573_/Q sky130_fd_sc_hd__dfrtp_1
X_1524_ _1524_/A VGND VGND VPWR VPWR _2435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1455_ _1455_/A VGND VGND VPWR VPWR _2475_/D sky130_fd_sc_hd__clkbuf_1
X_1386_ _1430_/A VGND VGND VPWR VPWR _1395_/S sky130_fd_sc_hd__clkbuf_2
X_2007_ _2011_/A VGND VGND VPWR VPWR _2007_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1240_ _2572_/Q _1233_/X _1234_/X _1239_/Y VGND VGND VPWR VPWR _2571_/D sky130_fd_sc_hd__a22o_1
X_1171_ _1171_/A _1171_/B VGND VGND VPWR VPWR _1172_/C sky130_fd_sc_hd__nor2_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput101 _2523_/Q VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__buf_2
X_2556_ _2560_/CLK _2556_/D _2313_/Y VGND VGND VPWR VPWR _2556_/Q sky130_fd_sc_hd__dfrtp_1
X_1507_ _1507_/A VGND VGND VPWR VPWR _2451_/D sky130_fd_sc_hd__clkbuf_1
X_2487_ _2487_/CLK _2487_/D _1980_/Y VGND VGND VPWR VPWR _2487_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1438_ _1438_/A VGND VGND VPWR VPWR _2482_/D sky130_fd_sc_hd__clkbuf_1
X_1369_ _2547_/Q _1194_/X _1364_/X _1368_/Y VGND VGND VPWR VPWR _2546_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2528_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput25 wbs_adr_i[30] VGND VGND VPWR VPWR _1171_/B sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_dat_i[10] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput14 wbs_adr_i[20] VGND VGND VPWR VPWR _1173_/B sky130_fd_sc_hd__clkbuf_1
Xinput47 wbs_dat_i[20] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 wbs_dat_i[30] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_2
X_2410_ _2549_/CLK _2410_/D _1885_/Y VGND VGND VPWR VPWR _2410_/Q sky130_fd_sc_hd__dfrtp_1
X_2341_ _2342_/A VGND VGND VPWR VPWR _2341_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2272_ _2272_/A _2477_/Q VGND VGND VPWR VPWR _2272_/Y sky130_fd_sc_hd__nand2_1
X_1223_ _2575_/Q _1209_/X _1220_/X _1222_/Y VGND VGND VPWR VPWR _2574_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1987_ _1987_/A VGND VGND VPWR VPWR _1987_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2539_ _2539_/CLK _2539_/D VGND VGND VPWR VPWR _2539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1912_/A VGND VGND VPWR VPWR _1910_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1841_ _1844_/A VGND VGND VPWR VPWR _1841_/Y sky130_fd_sc_hd__inv_2
X_1772_ _2585_/Q _2582_/Q _1771_/B VGND VGND VPWR VPWR _2585_/D sky130_fd_sc_hd__a21o_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2324_/A VGND VGND VPWR VPWR _2329_/A sky130_fd_sc_hd__buf_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _2245_/Y _2246_/X _2254_/Y VGND VGND VPWR VPWR _2539_/D sky130_fd_sc_hd__o21ai_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1206_ _2576_/Q VGND VGND VPWR VPWR _1206_/Y sky130_fd_sc_hd__inv_2
X_2186_ _2186_/A VGND VGND VPWR VPWR _2186_/X sky130_fd_sc_hd__buf_2
XFILLER_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2040_ _1361_/Y _2292_/B _2030_/X _2039_/Y VGND VGND VPWR VPWR _2040_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1824_ _2426_/Q VGND VGND VPWR VPWR _1828_/C sky130_fd_sc_hd__clkinv_2
X_1755_ _2581_/Q _2578_/Q VGND VGND VPWR VPWR _1755_/Y sky130_fd_sc_hd__nor2_1
X_1686_ _1777_/A _1686_/B _1686_/C _1686_/D VGND VGND VPWR VPWR _1687_/B sky130_fd_sc_hd__nor4_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2311_/A VGND VGND VPWR VPWR _2307_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2238_ _2238_/A VGND VGND VPWR VPWR _2272_/A sky130_fd_sc_hd__clkbuf_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2169_ _2530_/Q VGND VGND VPWR VPWR _2169_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1540_ _1540_/A VGND VGND VPWR VPWR _2428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1471_ _2467_/Q _2468_/Q _1473_/S VGND VGND VPWR VPWR _1472_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2023_ _2213_/A VGND VGND VPWR VPWR _2285_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ _1652_/C _2429_/Q _1805_/X _1806_/Y VGND VGND VPWR VPWR _1809_/A sky130_fd_sc_hd__o2bb2a_1
X_1738_ _1821_/C _2439_/Q _2405_/Q VGND VGND VPWR VPWR _2405_/D sky130_fd_sc_hd__a21o_1
X_1669_ _2385_/Q _2382_/Q VGND VGND VPWR VPWR _1673_/D sky130_fd_sc_hd__and2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2572_ _2575_/CLK _2572_/D _2333_/Y VGND VGND VPWR VPWR _2572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1523_ input54/X _2435_/Q _1523_/S VGND VGND VPWR VPWR _1524_/A sky130_fd_sc_hd__mux2_1
X_1454_ _2475_/Q _2476_/Q _1462_/S VGND VGND VPWR VPWR _1455_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1385_ _2448_/Q VGND VGND VPWR VPWR _1430_/A sky130_fd_sc_hd__buf_2
XFILLER_35_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2006_ _2006_/A VGND VGND VPWR VPWR _2011_/A sky130_fd_sc_hd__buf_2
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2403_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1170_ _2014_/A _1170_/B VGND VGND VPWR VPWR _1512_/A sky130_fd_sc_hd__nor2_4
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2555_ _2555_/CLK _2555_/D _2311_/Y VGND VGND VPWR VPWR _2555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1506_ _2451_/Q _2452_/Q _1506_/S VGND VGND VPWR VPWR _1507_/A sky130_fd_sc_hd__mux2_1
X_2486_ _2489_/CLK _2486_/D _1979_/Y VGND VGND VPWR VPWR _2486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1437_ _2482_/Q _2483_/Q _1439_/S VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__mux2_1
X_1368_ _1346_/X _2061_/B _1643_/A VGND VGND VPWR VPWR _1368_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1299_ _2559_/Q VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 wbs_adr_i[31] VGND VGND VPWR VPWR _1171_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 wbs_dat_i[11] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput15 wbs_adr_i[21] VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 wbs_dat_i[21] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 wbs_dat_i[31] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2340_ _2342_/A VGND VGND VPWR VPWR _2340_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2271_ _2285_/A _2285_/B _2436_/Q VGND VGND VPWR VPWR _2271_/Y sky130_fd_sc_hd__nor3b_1
X_1222_ _1212_/X _1214_/X _1221_/Y VGND VGND VPWR VPWR _1222_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1986_ _1987_/A VGND VGND VPWR VPWR _1986_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2538_ _2539_/CLK _2538_/D VGND VGND VPWR VPWR _2538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2469_ _2601_/CLK _2469_/D _1959_/Y VGND VGND VPWR VPWR _2469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ _1844_/A VGND VGND VPWR VPWR _1840_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1771_ _1771_/A _1771_/B VGND VGND VPWR VPWR _2584_/D sky130_fd_sc_hd__nor2_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2323_/A VGND VGND VPWR VPWR _2323_/Y sky130_fd_sc_hd__inv_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2248_/Y _2251_/Y _2253_/X VGND VGND VPWR VPWR _2254_/Y sky130_fd_sc_hd__o21ai_2
X_2185_ _2185_/A _2228_/B VGND VGND VPWR VPWR _2185_/Y sky130_fd_sc_hd__nor2_1
X_1205_ _2238_/A VGND VGND VPWR VPWR _2061_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1969_ _1975_/A VGND VGND VPWR VPWR _1974_/A sky130_fd_sc_hd__buf_4
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2578_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1823_ _2601_/Q _2598_/Q _1822_/B VGND VGND VPWR VPWR _2601_/D sky130_fd_sc_hd__a21o_1
X_1754_ _2581_/Q _2578_/Q VGND VGND VPWR VPWR _1754_/X sky130_fd_sc_hd__and2_1
X_1685_ _1631_/X _1686_/C _1686_/D _1686_/B VGND VGND VPWR VPWR _1687_/A sky130_fd_sc_hd__o22a_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2324_/A VGND VGND VPWR VPWR _2311_/A sky130_fd_sc_hd__buf_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2237_ _2237_/A VGND VGND VPWR VPWR _2237_/X sky130_fd_sc_hd__clkbuf_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2168_ _2159_/Y _2160_/X _2167_/Y VGND VGND VPWR VPWR _2529_/D sky130_fd_sc_hd__o21ai_1
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2099_ _2099_/A _2457_/Q VGND VGND VPWR VPWR _2099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1470_/A VGND VGND VPWR VPWR _2468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2022_ _2116_/A VGND VGND VPWR VPWR _2022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1806_ _2597_/Q _2594_/Q VGND VGND VPWR VPWR _1806_/Y sky130_fd_sc_hd__nor2_1
X_1737_ _1821_/C _2439_/Q _2405_/Q VGND VGND VPWR VPWR _1737_/X sky130_fd_sc_hd__and3_1
X_1668_ _2418_/Q VGND VGND VPWR VPWR _1673_/C sky130_fd_sc_hd__clkinv_2
X_1599_ _1599_/A VGND VGND VPWR VPWR _2442_/D sky130_fd_sc_hd__clkbuf_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2571_ _2577_/CLK _2571_/D _2332_/Y VGND VGND VPWR VPWR _2571_/Q sky130_fd_sc_hd__dfrtp_1
X_1522_ _1522_/A VGND VGND VPWR VPWR _2436_/D sky130_fd_sc_hd__clkbuf_1
X_1453_ _1486_/A VGND VGND VPWR VPWR _1462_/S sky130_fd_sc_hd__clkbuf_2
X_1384_ _1384_/A VGND VGND VPWR VPWR _2506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2005_ _2005_/A VGND VGND VPWR VPWR _2005_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2554_ _2555_/CLK _2554_/D _2310_/Y VGND VGND VPWR VPWR _2554_/Q sky130_fd_sc_hd__dfrtp_1
X_1505_ _1505_/A VGND VGND VPWR VPWR _2452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2485_ _2489_/CLK _2485_/D _1978_/Y VGND VGND VPWR VPWR _2485_/Q sky130_fd_sc_hd__dfrtp_1
X_1436_ _1436_/A VGND VGND VPWR VPWR _2483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1367_ _1672_/A VGND VGND VPWR VPWR _1643_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1298_ input39/X _1297_/X _1277_/X VGND VGND VPWR VPWR _1298_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 wbs_adr_i[3] VGND VGND VPWR VPWR _2013_/A sky130_fd_sc_hd__clkbuf_1
Xinput16 wbs_adr_i[22] VGND VGND VPWR VPWR _1174_/B sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_dat_i[12] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 wbs_dat_i[22] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2270_ _2542_/Q VGND VGND VPWR VPWR _2270_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1221_ _2574_/Q VGND VGND VPWR VPWR _1221_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1985_ _1987_/A VGND VGND VPWR VPWR _1985_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2537_ _2539_/CLK _2537_/D VGND VGND VPWR VPWR _2537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2468_ _2503_/CLK _2468_/D _1958_/Y VGND VGND VPWR VPWR _2468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1419_ _1430_/A VGND VGND VPWR VPWR _1428_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2399_ _2403_/CLK _2399_/D _1872_/Y VGND VGND VPWR VPWR _2399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ _1767_/X _1768_/Y _1789_/C _2435_/Q VGND VGND VPWR VPWR _1771_/B sky130_fd_sc_hd__and4bb_1
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _2323_/A VGND VGND VPWR VPWR _2322_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2253_ _2506_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2253_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2184_ _2532_/Q VGND VGND VPWR VPWR _2184_/Y sky130_fd_sc_hd__inv_2
X_1204_ _2026_/A VGND VGND VPWR VPWR _2238_/A sky130_fd_sc_hd__buf_4
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1968_ _1968_/A VGND VGND VPWR VPWR _1968_/Y sky130_fd_sc_hd__inv_2
X_1899_ _1900_/A VGND VGND VPWR VPWR _1899_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1822_ _1822_/A _1822_/B VGND VGND VPWR VPWR _2600_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1753_ _2579_/Q _2404_/Q _1752_/B VGND VGND VPWR VPWR _2579_/D sky130_fd_sc_hd__a21o_1
X_1684_ _2389_/Q _2386_/Q VGND VGND VPWR VPWR _1686_/B sky130_fd_sc_hd__nor2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2305_/A VGND VGND VPWR VPWR _2305_/Y sky130_fd_sc_hd__inv_2
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2264_/A _2236_/B _2432_/Q VGND VGND VPWR VPWR _2236_/Y sky130_fd_sc_hd__nor3b_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2167_ _2161_/Y _2164_/Y _2166_/X VGND VGND VPWR VPWR _2167_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_53_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2098_ _2098_/A _2161_/B VGND VGND VPWR VPWR _2098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2021_ _2146_/A VGND VGND VPWR VPWR _2116_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1805_ _2597_/Q _2594_/Q VGND VGND VPWR VPWR _1805_/X sky130_fd_sc_hd__and2_1
X_1736_ _2546_/Q VGND VGND VPWR VPWR _1821_/C sky130_fd_sc_hd__clkbuf_2
X_1667_ _2383_/Q _2380_/Q _1666_/B VGND VGND VPWR VPWR _2383_/D sky130_fd_sc_hd__a21o_1
X_1598_ _1596_/X _1614_/C _1598_/C VGND VGND VPWR VPWR _1599_/A sky130_fd_sc_hd__and3b_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2219_ _2212_/Y _2203_/X _2218_/Y VGND VGND VPWR VPWR _2535_/D sky130_fd_sc_hd__o21ai_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2570_ _2577_/CLK _2570_/D _2329_/Y VGND VGND VPWR VPWR _2570_/Q sky130_fd_sc_hd__dfrtp_1
X_1521_ input55/X _2436_/Q _1523_/S VGND VGND VPWR VPWR _1522_/A sky130_fd_sc_hd__mux2_1
X_1452_ _1452_/A VGND VGND VPWR VPWR _2476_/D sky130_fd_sc_hd__clkbuf_1
X_1383_ _2506_/Q _2507_/Q _1383_/S VGND VGND VPWR VPWR _1384_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2004_ _2005_/A VGND VGND VPWR VPWR _2004_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1719_ _1716_/X _1717_/Y _1751_/C _2411_/Q VGND VGND VPWR VPWR _1720_/B sky130_fd_sc_hd__and4bb_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2553_ _2553_/CLK _2553_/D _2309_/Y VGND VGND VPWR VPWR _2553_/Q sky130_fd_sc_hd__dfrtp_1
X_1504_ _2452_/Q _2453_/Q _1506_/S VGND VGND VPWR VPWR _1505_/A sky130_fd_sc_hd__mux2_1
X_2484_ _2484_/CLK _2484_/D _1977_/Y VGND VGND VPWR VPWR _2484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1435_ _2483_/Q _2484_/Q _1439_/S VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__mux2_1
X_1366_ _1722_/A VGND VGND VPWR VPWR _1672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1297_ _1297_/A VGND VGND VPWR VPWR _1297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2601_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput28 wbs_adr_i[4] VGND VGND VPWR VPWR _1167_/B sky130_fd_sc_hd__clkbuf_1
Xinput17 wbs_adr_i[23] VGND VGND VPWR VPWR _1174_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 wbs_dat_i[13] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1220_ input55/X _1219_/X _1339_/A VGND VGND VPWR VPWR _1220_/X sky130_fd_sc_hd__o21ba_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1984_ _1987_/A VGND VGND VPWR VPWR _1984_/Y sky130_fd_sc_hd__inv_2
X_2536_ _2536_/CLK _2536_/D VGND VGND VPWR VPWR _2536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2467_ _2497_/CLK _2467_/D _1956_/Y VGND VGND VPWR VPWR _2467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1418_ _1418_/A VGND VGND VPWR VPWR _2491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2398_ _2403_/CLK _2398_/D _1871_/Y VGND VGND VPWR VPWR _2398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1349_ _2551_/Q _1339_/X _1345_/X _1348_/Y VGND VGND VPWR VPWR _2550_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2323_/A VGND VGND VPWR VPWR _2321_/Y sky130_fd_sc_hd__inv_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2252_/A VGND VGND VPWR VPWR _2252_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1203_ _1512_/A _2028_/B _2028_/C VGND VGND VPWR VPWR _2026_/A sky130_fd_sc_hd__nand3_2
X_2183_ _2177_/Y _2160_/X _2182_/Y VGND VGND VPWR VPWR _2531_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1967_ _1968_/A VGND VGND VPWR VPWR _1967_/Y sky130_fd_sc_hd__inv_2
X_1898_ _1900_/A VGND VGND VPWR VPWR _1898_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2519_ _2520_/CLK _2519_/D VGND VGND VPWR VPWR _2519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2568_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ _1818_/X _1819_/Y _1821_/C _2427_/Q VGND VGND VPWR VPWR _1822_/B sky130_fd_sc_hd__and4bb_1
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1752_ _1752_/A _1752_/B VGND VGND VPWR VPWR _2578_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1683_ _2389_/Q _2386_/Q VGND VGND VPWR VPWR _1686_/D sky130_fd_sc_hd__and2_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2304_ _2305_/A VGND VGND VPWR VPWR _2304_/Y sky130_fd_sc_hd__inv_2
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2235_ _2538_/Q VGND VGND VPWR VPWR _2235_/Y sky130_fd_sc_hd__inv_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2166_ _2496_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2166_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2097_ _2522_/Q VGND VGND VPWR VPWR _2097_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2020_ _2231_/A VGND VGND VPWR VPWR _2146_/A sky130_fd_sc_hd__buf_2
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1804_ _2595_/Q _2592_/Q _1803_/B VGND VGND VPWR VPWR _2595_/D sky130_fd_sc_hd__a21o_1
X_1735_ _2403_/Q _2400_/Q _1734_/B VGND VGND VPWR VPWR _2403_/D sky130_fd_sc_hd__a21o_1
X_1666_ _1666_/A _1666_/B VGND VGND VPWR VPWR _2382_/D sky130_fd_sc_hd__nor2_1
X_1597_ _1588_/A _1593_/A _2442_/Q VGND VGND VPWR VPWR _1598_/C sky130_fd_sc_hd__a21o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2218_ _2214_/Y _2216_/Y _2217_/X VGND VGND VPWR VPWR _2218_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2149_ _2141_/Y _2116_/X _2148_/Y VGND VGND VPWR VPWR _2527_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1520_/A VGND VGND VPWR VPWR _2437_/D sky130_fd_sc_hd__clkbuf_1
X_1451_ _2476_/Q _2477_/Q _1451_/S VGND VGND VPWR VPWR _1452_/A sky130_fd_sc_hd__mux2_1
X_1382_ _1382_/A VGND VGND VPWR VPWR _2507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ _2005_/A VGND VGND VPWR VPWR _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1718_ _1702_/X _2411_/Q _1716_/X _1717_/Y VGND VGND VPWR VPWR _1720_/A sky130_fd_sc_hd__o2bb2a_1
X_1649_ _2379_/Q _2376_/Q VGND VGND VPWR VPWR _1649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2552_ _2553_/CLK _2552_/D _2308_/Y VGND VGND VPWR VPWR _2552_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _1503_/A VGND VGND VPWR VPWR _2453_/D sky130_fd_sc_hd__clkbuf_1
X_2483_ _2484_/CLK _2483_/D _1976_/Y VGND VGND VPWR VPWR _2483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1434_ _1434_/A VGND VGND VPWR VPWR _2484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1365_ _2546_/Q VGND VGND VPWR VPWR _1722_/A sky130_fd_sc_hd__inv_2
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1296_ _2561_/Q _1286_/X _1292_/X _1295_/Y VGND VGND VPWR VPWR _2560_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 wbs_adr_i[24] VGND VGND VPWR VPWR _1175_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput29 wbs_adr_i[5] VGND VGND VPWR VPWR _1167_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1983_ _1987_/A VGND VGND VPWR VPWR _1983_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2535_ _2568_/CLK _2535_/D VGND VGND VPWR VPWR _2535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2466_ _2497_/CLK _2466_/D _1955_/Y VGND VGND VPWR VPWR _2466_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1417_ _2491_/Q _2492_/Q _1417_/S VGND VGND VPWR VPWR _1418_/A sky130_fd_sc_hd__mux2_1
X_2397_ _2397_/CLK _2397_/D _1869_/Y VGND VGND VPWR VPWR _2397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1348_ _1346_/X _1341_/X _1347_/Y VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1279_ _2563_/Q VGND VGND VPWR VPWR _2178_/A sky130_fd_sc_hd__inv_2
XFILLER_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2323_/A VGND VGND VPWR VPWR _2320_/Y sky130_fd_sc_hd__inv_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2251_ _1238_/Y _2237_/X _2249_/X _2250_/Y VGND VGND VPWR VPWR _2251_/Y sky130_fd_sc_hd__o211ai_1
X_1202_ _2241_/A VGND VGND VPWR VPWR _1293_/A sky130_fd_sc_hd__buf_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2182_ _2178_/Y _2180_/Y _2181_/X VGND VGND VPWR VPWR _2182_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1966_ _1968_/A VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__inv_2
X_1897_ _1900_/A VGND VGND VPWR VPWR _1897_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2518_ _2520_/CLK _2518_/D VGND VGND VPWR VPWR _2518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2449_ _2484_/CLK _2449_/D _1934_/Y VGND VGND VPWR VPWR _2449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1820_ _1652_/C _2427_/Q _1818_/X _1819_/Y VGND VGND VPWR VPWR _1822_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1751_ _1748_/X _1749_/Y _1751_/C _2438_/Q VGND VGND VPWR VPWR _1752_/B sky130_fd_sc_hd__and4bb_1
X_1682_ _2416_/Q VGND VGND VPWR VPWR _1686_/C sky130_fd_sc_hd__inv_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2305_/A VGND VGND VPWR VPWR _2303_/Y sky130_fd_sc_hd__inv_2
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2227_/Y _2203_/X _2233_/Y VGND VGND VPWR VPWR _2537_/D sky130_fd_sc_hd__o21ai_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2165_/A VGND VGND VPWR VPWR _2165_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2096_ _2089_/Y _2071_/X _2095_/Y VGND VGND VPWR VPWR _2521_/D sky130_fd_sc_hd__o21ai_1
XFILLER_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1949_ _1949_/A VGND VGND VPWR VPWR _1949_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1803_ _1803_/A _1803_/B VGND VGND VPWR VPWR _2594_/D sky130_fd_sc_hd__nor2_1
X_1734_ _1734_/A _1734_/B VGND VGND VPWR VPWR _2402_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1665_ _1662_/X _1663_/Y _1706_/C _2419_/Q VGND VGND VPWR VPWR _1666_/B sky130_fd_sc_hd__and4bb_1
X_1596_ _2441_/Q _2440_/Q _2442_/Q VGND VGND VPWR VPWR _1596_/X sky130_fd_sc_hd__and3_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2502_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2217_/X sky130_fd_sc_hd__o31a_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ _2143_/Y _2145_/Y _2147_/X VGND VGND VPWR VPWR _2148_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2079_ _2486_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2079_/X sky130_fd_sc_hd__o31a_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1450_ _1450_/A VGND VGND VPWR VPWR _2477_/D sky130_fd_sc_hd__clkbuf_1
X_1381_ _2507_/Q _2508_/Q _1383_/S VGND VGND VPWR VPWR _1382_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2002_ _2005_/A VGND VGND VPWR VPWR _2002_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1717_ _2399_/Q _2396_/Q VGND VGND VPWR VPWR _1717_/Y sky130_fd_sc_hd__nor2_1
X_1648_ _2379_/Q _2376_/Q VGND VGND VPWR VPWR _1648_/X sky130_fd_sc_hd__and2_1
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A VGND VGND VPWR VPWR _2410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2551_ _2555_/CLK _2551_/D _2307_/Y VGND VGND VPWR VPWR _2551_/Q sky130_fd_sc_hd__dfrtp_1
X_1502_ _2453_/Q _2454_/Q _1506_/S VGND VGND VPWR VPWR _1503_/A sky130_fd_sc_hd__mux2_1
X_2482_ _2487_/CLK _2482_/D _1974_/Y VGND VGND VPWR VPWR _2482_/Q sky130_fd_sc_hd__dfrtp_2
X_1433_ _2484_/Q _2485_/Q _1439_/S VGND VGND VPWR VPWR _1434_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1364_ input35/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1364_/X sky130_fd_sc_hd__o21ba_1
X_1295_ _1293_/X _1288_/X _2151_/A VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2505_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 wbs_adr_i[25] VGND VGND VPWR VPWR _1175_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1982_ _2006_/A VGND VGND VPWR VPWR _1987_/A sky130_fd_sc_hd__buf_2
XFILLER_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2534_ _2536_/CLK _2534_/D VGND VGND VPWR VPWR _2534_/Q sky130_fd_sc_hd__dfxtp_1
X_2465_ _2465_/CLK _2465_/D _1954_/Y VGND VGND VPWR VPWR _2465_/Q sky130_fd_sc_hd__dfrtp_1
X_1416_ _1416_/A VGND VGND VPWR VPWR _2492_/D sky130_fd_sc_hd__clkbuf_1
X_2396_ _2397_/CLK _2396_/D _1868_/Y VGND VGND VPWR VPWR _2396_/Q sky130_fd_sc_hd__dfrtp_1
X_1347_ _2550_/Q VGND VGND VPWR VPWR _1347_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1278_ input43/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1278_/X sky130_fd_sc_hd__o21ba_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2250_ _2272_/A _2474_/Q VGND VGND VPWR VPWR _2250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1201_ _1512_/D VGND VGND VPWR VPWR _2241_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2181_ _2498_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2181_/X sky130_fd_sc_hd__o31a_1
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1965_ _1968_/A VGND VGND VPWR VPWR _1965_/Y sky130_fd_sc_hd__inv_2
X_1896_ _1900_/A VGND VGND VPWR VPWR _1896_/Y sky130_fd_sc_hd__inv_2
X_2517_ _2520_/CLK _2517_/D VGND VGND VPWR VPWR _2517_/Q sky130_fd_sc_hd__dfxtp_1
X_2448_ _2487_/CLK _2448_/D _1933_/Y VGND VGND VPWR VPWR _2448_/Q sky130_fd_sc_hd__dfrtp_4
X_2379_ _2447_/CLK _2379_/D _1847_/Y VGND VGND VPWR VPWR _2379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1750_ _1747_/X _2438_/Q _1748_/X _1749_/Y VGND VGND VPWR VPWR _1752_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1681_ _2387_/Q _2384_/Q _1680_/B VGND VGND VPWR VPWR _2387_/D sky130_fd_sc_hd__a21o_1
X_2302_ _2305_/A VGND VGND VPWR VPWR _2302_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2233_ _2228_/Y _2230_/Y _2232_/X VGND VGND VPWR VPWR _2233_/Y sky130_fd_sc_hd__o21ai_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _1636_/C _2118_/X _2162_/X _2163_/Y VGND VGND VPWR VPWR _2164_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2095_ _2091_/Y _2093_/Y _2094_/X VGND VGND VPWR VPWR _2095_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1948_ _1949_/A VGND VGND VPWR VPWR _1948_/Y sky130_fd_sc_hd__inv_2
X_1879_ _1881_/A VGND VGND VPWR VPWR _1879_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1802_ _1799_/X _1800_/Y _1821_/C _2430_/Q VGND VGND VPWR VPWR _1803_/B sky130_fd_sc_hd__and4bb_1
X_1733_ _1730_/X _1731_/Y _1751_/C _2409_/Q VGND VGND VPWR VPWR _1734_/B sky130_fd_sc_hd__and4bb_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1664_ _1647_/X _2419_/Q _1662_/X _1663_/Y VGND VGND VPWR VPWR _1666_/A sky130_fd_sc_hd__o2bb2a_1
X_1595_ _1588_/A _1593_/A _1594_/Y VGND VGND VPWR VPWR _2441_/D sky130_fd_sc_hd__a21oi_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2216_ _1258_/Y _2135_/X _2205_/X _2215_/Y VGND VGND VPWR VPWR _2216_/Y sky130_fd_sc_hd__o211ai_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2147_ _2494_/Q _2111_/X _2122_/X _2146_/X VGND VGND VPWR VPWR _2147_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2078_ _2165_/A VGND VGND VPWR VPWR _2078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1380_ _1380_/A VGND VGND VPWR VPWR _2508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2001_ _2005_/A VGND VGND VPWR VPWR _2001_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1716_ _2399_/Q _2396_/Q VGND VGND VPWR VPWR _1716_/X sky130_fd_sc_hd__and2_1
X_1647_ _1747_/A VGND VGND VPWR VPWR _1647_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ input57/X _2410_/Q _1578_/S VGND VGND VPWR VPWR _1579_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ _2550_/CLK _2550_/D _2305_/Y VGND VGND VPWR VPWR _2550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1501_ _1501_/A VGND VGND VPWR VPWR _2454_/D sky130_fd_sc_hd__clkbuf_1
X_2481_ _2487_/CLK _2481_/D _1973_/Y VGND VGND VPWR VPWR _2481_/Q sky130_fd_sc_hd__dfrtp_4
X_1432_ _1432_/A VGND VGND VPWR VPWR _2485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1363_ _2548_/Q _1339_/X _1360_/X _1362_/Y VGND VGND VPWR VPWR _2547_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1294_ _2560_/Q VGND VGND VPWR VPWR _2151_/A sky130_fd_sc_hd__inv_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1981_ input1/X VGND VGND VPWR VPWR _2006_/A sky130_fd_sc_hd__buf_2
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2533_ _2536_/CLK _2533_/D VGND VGND VPWR VPWR _2533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ _2465_/CLK _2464_/D _1953_/Y VGND VGND VPWR VPWR _2464_/Q sky130_fd_sc_hd__dfrtp_1
X_2395_ _2395_/CLK _2395_/D _1867_/Y VGND VGND VPWR VPWR _2395_/Q sky130_fd_sc_hd__dfrtp_1
X_1415_ _2492_/Q _2493_/Q _1417_/S VGND VGND VPWR VPWR _1416_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1346_ _1346_/A VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__clkbuf_2
X_1277_ _1374_/A VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _1200_/A VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__inv_2
X_2180_ _1621_/C _2118_/X _2162_/X _2179_/Y VGND VGND VPWR VPWR _2180_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1964_ _1968_/A VGND VGND VPWR VPWR _1964_/Y sky130_fd_sc_hd__inv_2
X_1895_ _1913_/A VGND VGND VPWR VPWR _1900_/A sky130_fd_sc_hd__buf_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2516_ _2549_/CLK _2516_/D VGND VGND VPWR VPWR _2516_/Q sky130_fd_sc_hd__dfxtp_1
X_2447_ _2447_/CLK _2447_/D _1931_/Y VGND VGND VPWR VPWR _2447_/Q sky130_fd_sc_hd__dfrtp_1
X_2378_ _2447_/CLK _2378_/D _1846_/Y VGND VGND VPWR VPWR _2378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ _2555_/Q _1311_/X _1326_/X _1328_/Y VGND VGND VPWR VPWR _2554_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1680_ _1680_/A _1680_/B VGND VGND VPWR VPWR _2386_/D sky130_fd_sc_hd__nor2_1
X_2301_ _2305_/A VGND VGND VPWR VPWR _2301_/Y sky130_fd_sc_hd__inv_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2232_ _2504_/Q _2198_/X _2208_/X _2231_/X VGND VGND VPWR VPWR _2232_/X sky130_fd_sc_hd__o31a_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2163_ _2187_/A _2464_/Q VGND VGND VPWR VPWR _2163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2094_ _2488_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2094_/X sky130_fd_sc_hd__o31a_1
XFILLER_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1947_ _1949_/A VGND VGND VPWR VPWR _1947_/Y sky130_fd_sc_hd__inv_2
X_1878_ _1881_/A VGND VGND VPWR VPWR _1878_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ _1652_/C _2430_/Q _1799_/X _1800_/Y VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__o2bb2a_1
X_1732_ _1702_/X _2409_/Q _1730_/X _1731_/Y VGND VGND VPWR VPWR _1734_/A sky130_fd_sc_hd__o2bb2a_1
X_1663_ _2383_/Q _2380_/Q VGND VGND VPWR VPWR _1663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1594_ _1588_/A _1593_/A _1194_/X VGND VGND VPWR VPWR _1594_/Y sky130_fd_sc_hd__o21ai_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _2229_/A _2470_/Q VGND VGND VPWR VPWR _2215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2146_ _2146_/A VGND VGND VPWR VPWR _2146_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2077_ _2252_/A VGND VGND VPWR VPWR _2165_/A sky130_fd_sc_hd__buf_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2593_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2000_ _2006_/A VGND VGND VPWR VPWR _2005_/A sky130_fd_sc_hd__buf_2
XFILLER_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1715_ _2397_/Q _2394_/Q _1714_/B VGND VGND VPWR VPWR _2397_/D sky130_fd_sc_hd__a21o_1
X_1646_ _2546_/Q VGND VGND VPWR VPWR _1747_/A sky130_fd_sc_hd__buf_2
X_1577_ _1577_/A VGND VGND VPWR VPWR _2411_/D sky130_fd_sc_hd__clkbuf_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2129_ _1308_/Y _2062_/X _2119_/X _2128_/Y VGND VGND VPWR VPWR _2129_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1500_ _2454_/Q _2455_/Q _1506_/S VGND VGND VPWR VPWR _1501_/A sky130_fd_sc_hd__mux2_1
X_2480_ _2504_/CLK _2480_/D _1972_/Y VGND VGND VPWR VPWR _2480_/Q sky130_fd_sc_hd__dfrtp_1
X_1431_ _2485_/Q _2486_/Q _1439_/S VGND VGND VPWR VPWR _1432_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput90 _2542_/Q VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__buf_2
X_1362_ _1346_/X _1341_/X _1361_/Y VGND VGND VPWR VPWR _1362_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1293_ _1293_/A VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1629_ _1629_/A _1629_/B VGND VGND VPWR VPWR _2372_/D sky130_fd_sc_hd__nor2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2567_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ _1980_/A VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2601_ _2601_/CLK _2601_/D _2367_/Y VGND VGND VPWR VPWR _2601_/Q sky130_fd_sc_hd__dfrtp_1
X_2532_ _2536_/CLK _2532_/D VGND VGND VPWR VPWR _2532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2463_ _2465_/CLK _2463_/D _1952_/Y VGND VGND VPWR VPWR _2463_/Q sky130_fd_sc_hd__dfrtp_1
X_2394_ _2397_/CLK _2394_/D _1866_/Y VGND VGND VPWR VPWR _2394_/Q sky130_fd_sc_hd__dfrtp_1
X_1414_ _1414_/A VGND VGND VPWR VPWR _2493_/D sky130_fd_sc_hd__clkbuf_1
X_1345_ input61/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1345_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1276_ _2565_/Q _1261_/X _1273_/X _1275_/Y VGND VGND VPWR VPWR _2564_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1963_ _1975_/A VGND VGND VPWR VPWR _1968_/A sky130_fd_sc_hd__buf_2
X_1894_ _1894_/A VGND VGND VPWR VPWR _1894_/Y sky130_fd_sc_hd__inv_2
X_2515_ _2549_/CLK _2515_/D VGND VGND VPWR VPWR _2515_/Q sky130_fd_sc_hd__dfxtp_1
X_2446_ _2446_/CLK _2446_/D _1930_/Y VGND VGND VPWR VPWR _2446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2377_ _2447_/CLK _2377_/D _1844_/Y VGND VGND VPWR VPWR _2377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1328_ _1320_/X _1313_/X _2098_/A VGND VGND VPWR VPWR _1328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1259_ _1242_/X _1237_/X _1258_/Y VGND VGND VPWR VPWR _1259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2300_ _2324_/A VGND VGND VPWR VPWR _2305_/A sky130_fd_sc_hd__buf_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2231_ _2231_/A VGND VGND VPWR VPWR _2231_/X sky130_fd_sc_hd__clkbuf_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2162_ _2249_/A VGND VGND VPWR VPWR _2162_/X sky130_fd_sc_hd__clkbuf_2
X_2093_ _1693_/C _1583_/S _2074_/X _2092_/Y VGND VGND VPWR VPWR _2093_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1946_ _1949_/A VGND VGND VPWR VPWR _1946_/Y sky130_fd_sc_hd__inv_2
X_1877_ _1881_/A VGND VGND VPWR VPWR _1877_/Y sky130_fd_sc_hd__inv_2
X_2429_ _2568_/CLK _2429_/D _1909_/Y VGND VGND VPWR VPWR _2429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ _2595_/Q _2592_/Q VGND VGND VPWR VPWR _1800_/Y sky130_fd_sc_hd__nor2_1
X_1731_ _2403_/Q _2400_/Q VGND VGND VPWR VPWR _1731_/Y sky130_fd_sc_hd__nor2_1
X_1662_ _2383_/Q _2380_/Q VGND VGND VPWR VPWR _1662_/X sky130_fd_sc_hd__and2_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1593_ _1593_/A _1593_/B VGND VGND VPWR VPWR _2440_/D sky130_fd_sc_hd__nor2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2264_/A _2236_/B _2429_/Q VGND VGND VPWR VPWR _2214_/Y sky130_fd_sc_hd__nor3b_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _1299_/Y _2135_/X _2119_/X _2144_/Y VGND VGND VPWR VPWR _2145_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ _1342_/Y _2062_/X _2074_/X _2075_/Y VGND VGND VPWR VPWR _2076_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ _1931_/A VGND VGND VPWR VPWR _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1714_ _1714_/A _1714_/B VGND VGND VPWR VPWR _2396_/D sky130_fd_sc_hd__nor2_1
X_1645_ _2377_/Q _2374_/Q _1644_/B VGND VGND VPWR VPWR _2377_/D sky130_fd_sc_hd__a21o_1
X_1576_ input60/X _2411_/Q _1578_/S VGND VGND VPWR VPWR _1577_/A sky130_fd_sc_hd__mux2_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2128_ _2144_/A _2460_/Q VGND VGND VPWR VPWR _2128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2059_ _2052_/Y _2022_/X _2058_/Y VGND VGND VPWR VPWR _2517_/D sky130_fd_sc_hd__o21ai_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A VGND VGND VPWR VPWR _1439_/S sky130_fd_sc_hd__buf_2
X_1361_ _2547_/Q VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput80 _2533_/Q VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput91 _2543_/Q VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_1292_ input40/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2492_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1628_ _1643_/A _1628_/B _1628_/C _1628_/D VGND VGND VPWR VPWR _1629_/B sky130_fd_sc_hd__nor4_1
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1559_ input37/X _2419_/Q _1567_/S VGND VGND VPWR VPWR _1560_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2600_ _2601_/CLK _2600_/D _2366_/Y VGND VGND VPWR VPWR _2600_/Q sky130_fd_sc_hd__dfrtp_1
X_2531_ _2536_/CLK _2531_/D VGND VGND VPWR VPWR _2531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2462_ _2465_/CLK _2462_/D _1949_/Y VGND VGND VPWR VPWR _2462_/Q sky130_fd_sc_hd__dfrtp_1
X_2393_ _2395_/CLK _2393_/D _1865_/Y VGND VGND VPWR VPWR _2393_/Q sky130_fd_sc_hd__dfrtp_1
X_1413_ _2493_/Q _2494_/Q _1417_/S VGND VGND VPWR VPWR _1414_/A sky130_fd_sc_hd__mux2_1
X_1344_ _2552_/Q _1339_/X _1340_/X _1343_/Y VGND VGND VPWR VPWR _2551_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1275_ _1268_/X _1263_/X _2185_/A VGND VGND VPWR VPWR _1275_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _1962_/A VGND VGND VPWR VPWR _1962_/Y sky130_fd_sc_hd__inv_2
X_1893_ _1894_/A VGND VGND VPWR VPWR _1893_/Y sky130_fd_sc_hd__inv_2
X_2514_ _2549_/CLK _2514_/D VGND VGND VPWR VPWR _2514_/Q sky130_fd_sc_hd__dfxtp_1
X_2445_ _2446_/CLK _2445_/D _1929_/Y VGND VGND VPWR VPWR _2445_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ _2447_/CLK _2376_/D _1843_/Y VGND VGND VPWR VPWR _2376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1327_ _2554_/Q VGND VGND VPWR VPWR _2098_/A sky130_fd_sc_hd__inv_2
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1258_ _2567_/Q VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1189_ _2213_/A _1512_/A _2028_/B _2028_/C VGND VGND VPWR VPWR _1324_/A sky130_fd_sc_hd__nand4_1
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _1796_/C _2186_/X _2205_/X _2229_/Y VGND VGND VPWR VPWR _2230_/Y sky130_fd_sc_hd__o211ai_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ _2161_/A _2161_/B VGND VGND VPWR VPWR _2161_/Y sky130_fd_sc_hd__nor2_1
X_2092_ _2099_/A _2456_/Q VGND VGND VPWR VPWR _2092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1945_ _1949_/A VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1876_ _1882_/A VGND VGND VPWR VPWR _1881_/A sky130_fd_sc_hd__buf_4
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2428_ _2536_/CLK _2428_/D _1908_/Y VGND VGND VPWR VPWR _2428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2359_ _2360_/A VGND VGND VPWR VPWR _2359_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1730_ _2403_/Q _2400_/Q VGND VGND VPWR VPWR _1730_/X sky130_fd_sc_hd__and2_1
X_1661_ _2381_/Q _2378_/Q _1660_/B VGND VGND VPWR VPWR _2381_/D sky130_fd_sc_hd__a21o_1
X_1592_ _2440_/Q VGND VGND VPWR VPWR _1593_/A sky130_fd_sc_hd__clkbuf_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2213_ _2213_/A VGND VGND VPWR VPWR _2264_/A sky130_fd_sc_hd__clkbuf_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2144_ _2144_/A _2462_/Q VGND VGND VPWR VPWR _2144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2075_ _2099_/A _2454_/Q VGND VGND VPWR VPWR _2075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1928_ _1931_/A VGND VGND VPWR VPWR _1928_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ _1863_/A VGND VGND VPWR VPWR _1859_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_2_0_wb_clk_i/X VGND VGND VPWR VPWR _2575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1713_ _1709_/X _1710_/Y _1751_/C _2412_/Q VGND VGND VPWR VPWR _1714_/B sky130_fd_sc_hd__and4bb_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_0 _2034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1644_ _1644_/A _1644_/B VGND VGND VPWR VPWR _2376_/D sky130_fd_sc_hd__nor2_1
X_1575_ _1575_/A VGND VGND VPWR VPWR _2412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _2194_/A _2134_/B _2419_/Q VGND VGND VPWR VPWR _2127_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2058_ _2053_/Y _2055_/Y _2057_/X VGND VGND VPWR VPWR _2058_/Y sky130_fd_sc_hd__o21ai_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput70 _2514_/Q VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__buf_2
X_1360_ input46/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1360_/X sky130_fd_sc_hd__o21ba_1
Xoutput92 _2516_/Q VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput81 _2515_/Q VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _2562_/Q _1286_/X _1287_/X _1290_/Y VGND VGND VPWR VPWR _2561_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1627_ _1828_/A _1628_/C _1628_/D _1628_/B VGND VGND VPWR VPWR _1629_/A sky130_fd_sc_hd__o22a_1
X_1558_ _1558_/A VGND VGND VPWR VPWR _1567_/S sky130_fd_sc_hd__buf_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1489_ _2459_/Q _2460_/Q _1495_/S VGND VGND VPWR VPWR _1490_/A sky130_fd_sc_hd__mux2_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2550_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2530_ _2536_/CLK _2530_/D VGND VGND VPWR VPWR _2530_/Q sky130_fd_sc_hd__dfxtp_1
X_2461_ _2495_/CLK _2461_/D _1948_/Y VGND VGND VPWR VPWR _2461_/Q sky130_fd_sc_hd__dfrtp_1
X_1412_ _1412_/A VGND VGND VPWR VPWR _2494_/D sky130_fd_sc_hd__clkbuf_1
X_2392_ _2395_/CLK _2392_/D _1863_/Y VGND VGND VPWR VPWR _2392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1343_ _1320_/X _1341_/X _1342_/Y VGND VGND VPWR VPWR _1343_/Y sky130_fd_sc_hd__o21ai_1
X_1274_ _2564_/Q VGND VGND VPWR VPWR _2185_/A sky130_fd_sc_hd__inv_2
XFILLER_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1961_ _1962_/A VGND VGND VPWR VPWR _1961_/Y sky130_fd_sc_hd__inv_2
X_1892_ _1894_/A VGND VGND VPWR VPWR _1892_/Y sky130_fd_sc_hd__inv_2
X_2513_ _2550_/CLK _2513_/D VGND VGND VPWR VPWR _2513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2444_ _2446_/CLK _2444_/D _1928_/Y VGND VGND VPWR VPWR _2444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2375_ _2406_/CLK _2375_/D _1842_/Y VGND VGND VPWR VPWR _2375_/Q sky130_fd_sc_hd__dfrtp_1
X_1326_ input65/X _1325_/X _1302_/X VGND VGND VPWR VPWR _1326_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1257_ input48/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__o21ba_1
X_1188_ _1188_/A _1188_/B VGND VGND VPWR VPWR _2028_/C sky130_fd_sc_hd__nor2_4
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2246_/A VGND VGND VPWR VPWR _2160_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ _2091_/A _2161_/B VGND VGND VPWR VPWR _2091_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1944_ _1944_/A VGND VGND VPWR VPWR _1949_/A sky130_fd_sc_hd__buf_2
X_1875_ _1875_/A VGND VGND VPWR VPWR _1875_/Y sky130_fd_sc_hd__inv_2
X_2427_ _2536_/CLK _2427_/D _1906_/Y VGND VGND VPWR VPWR _2427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2358_ _2360_/A VGND VGND VPWR VPWR _2358_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1309_ _1293_/X _1288_/X _1308_/Y VGND VGND VPWR VPWR _1309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2289_ _2285_/Y _2287_/Y _2288_/X VGND VGND VPWR VPWR _2289_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1660_ _1660_/A _1660_/B VGND VGND VPWR VPWR _2380_/D sky130_fd_sc_hd__nor2_1
X_1591_ _1194_/X _1191_/X _1593_/B VGND VGND VPWR VPWR _2448_/D sky130_fd_sc_hd__o21ai_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2535_/Q VGND VGND VPWR VPWR _2212_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2143_ _2194_/A _2236_/B _2421_/Q VGND VGND VPWR VPWR _2143_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2074_ _2074_/A VGND VGND VPWR VPWR _2074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1927_ _1931_/A VGND VGND VPWR VPWR _1927_/Y sky130_fd_sc_hd__inv_2
X_1858_ _1882_/A VGND VGND VPWR VPWR _1863_/A sky130_fd_sc_hd__buf_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1789_ _1786_/X _1787_/Y _1789_/C _2432_/Q VGND VGND VPWR VPWR _1790_/B sky130_fd_sc_hd__and4bb_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1712_ _1747_/A VGND VGND VPWR VPWR _1751_/C sky130_fd_sc_hd__buf_4
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 _2448_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ _1643_/A _1643_/B _1643_/C _1643_/D VGND VGND VPWR VPWR _1644_/B sky130_fd_sc_hd__nor4_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1574_ input61/X _2412_/Q _1578_/S VGND VGND VPWR VPWR _1575_/A sky130_fd_sc_hd__mux2_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2126_ _2525_/Q VGND VGND VPWR VPWR _2126_/Y sky130_fd_sc_hd__inv_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2057_ _2484_/Q _1346_/A _2016_/X _2056_/X VGND VGND VPWR VPWR _2057_/X sky130_fd_sc_hd__o31a_1
XFILLER_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput93 _2544_/Q VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput71 _2524_/Q VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput82 _2534_/Q VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_1290_ _1268_/X _1288_/X _2161_/A VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _2373_/Q _2370_/Q VGND VGND VPWR VPWR _1628_/B sky130_fd_sc_hd__nor2_1
X_1557_ _1557_/A VGND VGND VPWR VPWR _2420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1488_ _1488_/A VGND VGND VPWR VPWR _2460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ _2144_/A _2458_/Q VGND VGND VPWR VPWR _2109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2447_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ _2487_/CLK _2460_/D _1947_/Y VGND VGND VPWR VPWR _2460_/Q sky130_fd_sc_hd__dfrtp_1
X_1411_ _2494_/Q _2495_/Q _1417_/S VGND VGND VPWR VPWR _1412_/A sky130_fd_sc_hd__mux2_1
X_2391_ _2397_/CLK _2391_/D _1862_/Y VGND VGND VPWR VPWR _2391_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1342_ _2551_/Q VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1273_ input44/X _1272_/X _1252_/X VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__o21ba_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2589_ _2589_/CLK _2589_/D _2353_/Y VGND VGND VPWR VPWR _2589_/Q sky130_fd_sc_hd__dfrtp_1
X_1609_ _1609_/A VGND VGND VPWR VPWR _2445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ _1962_/A VGND VGND VPWR VPWR _1960_/Y sky130_fd_sc_hd__inv_2
X_1891_ _1894_/A VGND VGND VPWR VPWR _1891_/Y sky130_fd_sc_hd__inv_2
X_2512_ _2578_/CLK _2512_/D _2011_/Y VGND VGND VPWR VPWR _2512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2443_ _2446_/CLK _2443_/D _1927_/Y VGND VGND VPWR VPWR _2443_/Q sky130_fd_sc_hd__dfrtp_1
X_2374_ _2465_/CLK _2374_/D _1841_/Y VGND VGND VPWR VPWR _2374_/Q sky130_fd_sc_hd__dfrtp_1
X_1325_ _2170_/A VGND VGND VPWR VPWR _1325_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1256_ _2569_/Q _1233_/X _1253_/X _1255_/Y VGND VGND VPWR VPWR _2568_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1187_ _1187_/A _1187_/B _1187_/C _1187_/D VGND VGND VPWR VPWR _1188_/B sky130_fd_sc_hd__nand4_1
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2090_ _2170_/A VGND VGND VPWR VPWR _2161_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1943_ _1943_/A VGND VGND VPWR VPWR _1943_/Y sky130_fd_sc_hd__inv_2
X_1874_ _1875_/A VGND VGND VPWR VPWR _1874_/Y sky130_fd_sc_hd__inv_2
X_2426_ _2567_/CLK _2426_/D _1905_/Y VGND VGND VPWR VPWR _2426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2357_ _2360_/A VGND VGND VPWR VPWR _2357_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1308_ _2557_/Q VGND VGND VPWR VPWR _1308_/Y sky130_fd_sc_hd__inv_2
X_2288_ _2511_/Q _2066_/A _2165_/A _2032_/X VGND VGND VPWR VPWR _2288_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1239_ _1212_/X _1237_/X _1238_/Y VGND VGND VPWR VPWR _1239_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1590_ _1586_/X _1588_/X _1614_/C VGND VGND VPWR VPWR _1593_/B sky130_fd_sc_hd__o21ai_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2202_/Y _2203_/X _2210_/Y VGND VGND VPWR VPWR _2534_/D sky130_fd_sc_hd__o21ai_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2142_ _2247_/A VGND VGND VPWR VPWR _2236_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2073_ _2083_/A _2134_/B _2413_/Q VGND VGND VPWR VPWR _2073_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1926_ _1944_/A VGND VGND VPWR VPWR _1931_/A sky130_fd_sc_hd__buf_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1857_ _2361_/A VGND VGND VPWR VPWR _1882_/A sky130_fd_sc_hd__buf_2
X_1788_ _1652_/C _2432_/Q _1786_/X _1787_/Y VGND VGND VPWR VPWR _1790_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2409_ _2453_/CLK _2409_/D _1884_/Y VGND VGND VPWR VPWR _2409_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2561_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1711_ _1702_/X _2412_/Q _1709_/X _1710_/Y VGND VGND VPWR VPWR _1714_/A sky130_fd_sc_hd__o2bb2a_1
XANTENNA_2 _2406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _1631_/X _1643_/C _1643_/D _1643_/B VGND VGND VPWR VPWR _1644_/A sky130_fd_sc_hd__o22a_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1573_ _1573_/A VGND VGND VPWR VPWR _2413_/D sky130_fd_sc_hd__clkbuf_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _2115_/Y _2116_/X _2124_/Y VGND VGND VPWR VPWR _2524_/D sky130_fd_sc_hd__o21ai_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2056_ _2146_/A VGND VGND VPWR VPWR _2056_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1909_ _1912_/A VGND VGND VPWR VPWR _1909_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput94 _2545_/Q VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput72 _2525_/Q VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput83 _2535_/Q VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1625_ _2373_/Q _2370_/Q VGND VGND VPWR VPWR _1628_/D sky130_fd_sc_hd__and2_1
X_1556_ input38/X _2420_/Q _1556_/S VGND VGND VPWR VPWR _1557_/A sky130_fd_sc_hd__mux2_1
X_1487_ _2460_/Q _2461_/Q _1495_/S VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__mux2_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2108_ _2247_/A VGND VGND VPWR VPWR _2144_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2039_ _2054_/A _2450_/Q VGND VGND VPWR VPWR _2039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1410_ _1410_/A VGND VGND VPWR VPWR _2495_/D sky130_fd_sc_hd__clkbuf_1
X_2390_ _2395_/CLK _2390_/D _1861_/Y VGND VGND VPWR VPWR _2390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1341_ _2054_/A VGND VGND VPWR VPWR _1341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1272_ _1297_/A VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1608_ _1612_/C _1608_/B _1608_/C VGND VGND VPWR VPWR _1609_/A sky130_fd_sc_hd__and3b_1
X_2588_ _2589_/CLK _2588_/D _2352_/Y VGND VGND VPWR VPWR _2588_/Q sky130_fd_sc_hd__dfrtp_1
X_1539_ input47/X _2428_/Q _1545_/S VGND VGND VPWR VPWR _1540_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1890_ _1894_/A VGND VGND VPWR VPWR _1890_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ _2578_/CLK _2511_/D _2010_/Y VGND VGND VPWR VPWR _2511_/Q sky130_fd_sc_hd__dfrtp_1
X_2442_ _2597_/CLK _2442_/D _1925_/Y VGND VGND VPWR VPWR _2442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2373_ _2447_/CLK _2373_/D _1840_/Y VGND VGND VPWR VPWR _2373_/Q sky130_fd_sc_hd__dfrtp_1
X_1324_ _1324_/A VGND VGND VPWR VPWR _2170_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1255_ _1242_/X _1237_/X _1254_/Y VGND VGND VPWR VPWR _1255_/Y sky130_fd_sc_hd__o21ai_1
X_1186_ input8/X input7/X VGND VGND VPWR VPWR _1187_/D sky130_fd_sc_hd__nor2_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1942_ _1943_/A VGND VGND VPWR VPWR _1942_/Y sky130_fd_sc_hd__inv_2
X_1873_ _1875_/A VGND VGND VPWR VPWR _1873_/Y sky130_fd_sc_hd__inv_2
X_2425_ _2529_/CLK _2425_/D _1904_/Y VGND VGND VPWR VPWR _2425_/Q sky130_fd_sc_hd__dfrtp_1
X_2356_ _2360_/A VGND VGND VPWR VPWR _2356_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1307_ input37/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__o21ba_1
X_2287_ _1206_/Y _1297_/A _2074_/A _2286_/Y VGND VGND VPWR VPWR _2287_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1238_ _2571_/Q VGND VGND VPWR VPWR _1238_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1169_ _2013_/A _2012_/B VGND VGND VPWR VPWR _1170_/B sky130_fd_sc_hd__or2b_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2210_ _2204_/Y _2207_/Y _2209_/X VGND VGND VPWR VPWR _2210_/Y sky130_fd_sc_hd__o21ai_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2141_ _2527_/Q VGND VGND VPWR VPWR _2141_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2072_ _2294_/A VGND VGND VPWR VPWR _2134_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1925_ _1925_/A VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_2_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2484_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1856_ _1856_/A VGND VGND VPWR VPWR _1856_/Y sky130_fd_sc_hd__inv_2
X_1787_ _2591_/Q _2588_/Q VGND VGND VPWR VPWR _1787_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2408_ _2453_/CLK _2408_/D _1883_/Y VGND VGND VPWR VPWR _2408_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2339_ _2342_/A VGND VGND VPWR VPWR _2339_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1710_ _2397_/Q _2394_/Q VGND VGND VPWR VPWR _1710_/Y sky130_fd_sc_hd__nor2_1
X_1641_ _2377_/Q _2374_/Q VGND VGND VPWR VPWR _1643_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1572_ input62/X _2413_/Q _1578_/S VGND VGND VPWR VPWR _1573_/A sky130_fd_sc_hd__mux2_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2124_ _2117_/Y _2121_/Y _2123_/X VGND VGND VPWR VPWR _2124_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2055_ _1352_/Y _2292_/B _2030_/X _2054_/Y VGND VGND VPWR VPWR _2055_/Y sky130_fd_sc_hd__o211ai_1
X_1908_ _1912_/A VGND VGND VPWR VPWR _1908_/Y sky130_fd_sc_hd__inv_2
X_1839_ _2367_/A VGND VGND VPWR VPWR _1844_/A sky130_fd_sc_hd__buf_2
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput73 _2526_/Q VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput84 _2536_/Q VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput95 _2517_/Q VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1624_ _2424_/Q VGND VGND VPWR VPWR _1628_/C sky130_fd_sc_hd__clkinv_2
X_1555_ _1555_/A VGND VGND VPWR VPWR _2421_/D sky130_fd_sc_hd__clkbuf_1
X_1486_ _1486_/A VGND VGND VPWR VPWR _1495_/S sky130_fd_sc_hd__buf_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2107_ _2194_/A _2134_/B _2417_/Q VGND VGND VPWR VPWR _2107_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2038_ _2083_/A _2061_/B _2409_/Q VGND VGND VPWR VPWR _2038_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ input62/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3_0_wb_clk_i/X VGND VGND VPWR VPWR _2587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1271_ _2566_/Q _1261_/X _1267_/X _1270_/Y VGND VGND VPWR VPWR _2565_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1607_ _2443_/Q _1586_/B _1596_/X _2445_/Q VGND VGND VPWR VPWR _1608_/C sky130_fd_sc_hd__a31o_1
X_2587_ _2587_/CLK _2587_/D _2351_/Y VGND VGND VPWR VPWR _2587_/Q sky130_fd_sc_hd__dfrtp_1
X_1538_ _1538_/A VGND VGND VPWR VPWR _2429_/D sky130_fd_sc_hd__clkbuf_1
X_1469_ _2468_/Q _2469_/Q _1473_/S VGND VGND VPWR VPWR _1470_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2510_ _2510_/CLK _2510_/D _2009_/Y VGND VGND VPWR VPWR _2510_/Q sky130_fd_sc_hd__dfrtp_1
X_2441_ _2597_/CLK _2441_/D _1924_/Y VGND VGND VPWR VPWR _2441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2372_ _2497_/CLK _2372_/D _1838_/Y VGND VGND VPWR VPWR _2372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1323_ _2556_/Q _1311_/X _1317_/X _1322_/Y VGND VGND VPWR VPWR _2555_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1254_ _2568_/Q VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1185_ input6/X input5/X VGND VGND VPWR VPWR _1187_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1941_ _1943_/A VGND VGND VPWR VPWR _1941_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ _1875_/A VGND VGND VPWR VPWR _1872_/Y sky130_fd_sc_hd__inv_2
X_2424_ _2529_/CLK _2424_/D _1903_/Y VGND VGND VPWR VPWR _2424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2355_ _2355_/A VGND VGND VPWR VPWR _2360_/A sky130_fd_sc_hd__buf_2
XFILLER_69_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1306_ _2559_/Q _1286_/X _1303_/X _1305_/Y VGND VGND VPWR VPWR _2558_/D sky130_fd_sc_hd__a22o_1
X_2286_ _2294_/A _2479_/Q VGND VGND VPWR VPWR _2286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1237_ _2024_/B VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1168_ _1165_/Y _1168_/B _1168_/C VGND VGND VPWR VPWR _2014_/A sky130_fd_sc_hd__nand3b_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2133_/Y _2116_/X _2139_/Y VGND VGND VPWR VPWR _2526_/D sky130_fd_sc_hd__o21ai_1
X_2071_ _2116_/A VGND VGND VPWR VPWR _2071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1924_ _1925_/A VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1855_ _1856_/A VGND VGND VPWR VPWR _1855_/Y sky130_fd_sc_hd__inv_2
X_1786_ _2591_/Q _2588_/Q VGND VGND VPWR VPWR _1786_/X sky130_fd_sc_hd__and2_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2407_ _2487_/CLK _2407_/D _1881_/Y VGND VGND VPWR VPWR _2407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2338_ _2342_/A VGND VGND VPWR VPWR _2338_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2269_ _2263_/Y _2246_/X _2268_/Y VGND VGND VPWR VPWR _2541_/D sky130_fd_sc_hd__o21ai_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1640_ _2377_/Q _2374_/Q VGND VGND VPWR VPWR _1643_/D sky130_fd_sc_hd__and2_1
X_1571_ _1571_/A VGND VGND VPWR VPWR _2414_/D sky130_fd_sc_hd__clkbuf_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ _2491_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2123_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2054_ _2054_/A _2452_/Q VGND VGND VPWR VPWR _2054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1907_ _1913_/A VGND VGND VPWR VPWR _1912_/A sky130_fd_sc_hd__buf_2
X_1838_ _1838_/A VGND VGND VPWR VPWR _1838_/Y sky130_fd_sc_hd__inv_2
X_1769_ _1747_/X _2435_/Q _1767_/X _1768_/Y VGND VGND VPWR VPWR _1771_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput74 _2527_/Q VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput85 _2537_/Q VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput96 _2518_/Q VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1623_ _2371_/Q _2368_/Q _1622_/B VGND VGND VPWR VPWR _2371_/D sky130_fd_sc_hd__a21o_1
X_1554_ input39/X _2421_/Q _1556_/S VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__mux2_1
X_1485_ _1485_/A VGND VGND VPWR VPWR _2461_/D sky130_fd_sc_hd__clkbuf_1
.ends

