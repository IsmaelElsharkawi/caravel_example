magic
tech sky130A
magscale 1 2
timestamp 1650980003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 8 179202 117552
<< metal2 >>
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9310 0 9366 800
rect 10966 0 11022 800
rect 12714 0 12770 800
rect 14370 0 14426 800
rect 16118 0 16174 800
rect 17774 0 17830 800
rect 19522 0 19578 800
rect 21178 0 21234 800
rect 22926 0 22982 800
rect 24582 0 24638 800
rect 26238 0 26294 800
rect 27986 0 28042 800
rect 29642 0 29698 800
rect 31390 0 31446 800
rect 33046 0 33102 800
rect 34794 0 34850 800
rect 36450 0 36506 800
rect 38198 0 38254 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 45006 0 45062 800
rect 46662 0 46718 800
rect 48318 0 48374 800
rect 50066 0 50122 800
rect 51722 0 51778 800
rect 53470 0 53526 800
rect 55126 0 55182 800
rect 56874 0 56930 800
rect 58530 0 58586 800
rect 60278 0 60334 800
rect 61934 0 61990 800
rect 63682 0 63738 800
rect 65338 0 65394 800
rect 67086 0 67142 800
rect 68742 0 68798 800
rect 70398 0 70454 800
rect 72146 0 72202 800
rect 73802 0 73858 800
rect 75550 0 75606 800
rect 77206 0 77262 800
rect 78954 0 79010 800
rect 80610 0 80666 800
rect 82358 0 82414 800
rect 84014 0 84070 800
rect 85762 0 85818 800
rect 87418 0 87474 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94226 0 94282 800
rect 95882 0 95938 800
rect 97630 0 97686 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102690 0 102746 800
rect 104438 0 104494 800
rect 106094 0 106150 800
rect 107842 0 107898 800
rect 109498 0 109554 800
rect 111246 0 111302 800
rect 112902 0 112958 800
rect 114558 0 114614 800
rect 116306 0 116362 800
rect 117962 0 118018 800
rect 119710 0 119766 800
rect 121366 0 121422 800
rect 123114 0 123170 800
rect 124770 0 124826 800
rect 126518 0 126574 800
rect 128174 0 128230 800
rect 129922 0 129978 800
rect 131578 0 131634 800
rect 133326 0 133382 800
rect 134982 0 135038 800
rect 136638 0 136694 800
rect 138386 0 138442 800
rect 140042 0 140098 800
rect 141790 0 141846 800
rect 143446 0 143502 800
rect 145194 0 145250 800
rect 146850 0 146906 800
rect 148598 0 148654 800
rect 150254 0 150310 800
rect 152002 0 152058 800
rect 153658 0 153714 800
rect 155406 0 155462 800
rect 157062 0 157118 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162122 0 162178 800
rect 163870 0 163926 800
rect 165526 0 165582 800
rect 167274 0 167330 800
rect 168930 0 168986 800
rect 170678 0 170734 800
rect 172334 0 172390 800
rect 174082 0 174138 800
rect 175738 0 175794 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 846 856 179196 117552
rect 958 2 2446 856
rect 2614 2 4102 856
rect 4270 2 5850 856
rect 6018 2 7506 856
rect 7674 2 9254 856
rect 9422 2 10910 856
rect 11078 2 12658 856
rect 12826 2 14314 856
rect 14482 2 16062 856
rect 16230 2 17718 856
rect 17886 2 19466 856
rect 19634 2 21122 856
rect 21290 2 22870 856
rect 23038 2 24526 856
rect 24694 2 26182 856
rect 26350 2 27930 856
rect 28098 2 29586 856
rect 29754 2 31334 856
rect 31502 2 32990 856
rect 33158 2 34738 856
rect 34906 2 36394 856
rect 36562 2 38142 856
rect 38310 2 39798 856
rect 39966 2 41546 856
rect 41714 2 43202 856
rect 43370 2 44950 856
rect 45118 2 46606 856
rect 46774 2 48262 856
rect 48430 2 50010 856
rect 50178 2 51666 856
rect 51834 2 53414 856
rect 53582 2 55070 856
rect 55238 2 56818 856
rect 56986 2 58474 856
rect 58642 2 60222 856
rect 60390 2 61878 856
rect 62046 2 63626 856
rect 63794 2 65282 856
rect 65450 2 67030 856
rect 67198 2 68686 856
rect 68854 2 70342 856
rect 70510 2 72090 856
rect 72258 2 73746 856
rect 73914 2 75494 856
rect 75662 2 77150 856
rect 77318 2 78898 856
rect 79066 2 80554 856
rect 80722 2 82302 856
rect 82470 2 83958 856
rect 84126 2 85706 856
rect 85874 2 87362 856
rect 87530 2 89110 856
rect 89278 2 90766 856
rect 90934 2 92422 856
rect 92590 2 94170 856
rect 94338 2 95826 856
rect 95994 2 97574 856
rect 97742 2 99230 856
rect 99398 2 100978 856
rect 101146 2 102634 856
rect 102802 2 104382 856
rect 104550 2 106038 856
rect 106206 2 107786 856
rect 107954 2 109442 856
rect 109610 2 111190 856
rect 111358 2 112846 856
rect 113014 2 114502 856
rect 114670 2 116250 856
rect 116418 2 117906 856
rect 118074 2 119654 856
rect 119822 2 121310 856
rect 121478 2 123058 856
rect 123226 2 124714 856
rect 124882 2 126462 856
rect 126630 2 128118 856
rect 128286 2 129866 856
rect 130034 2 131522 856
rect 131690 2 133270 856
rect 133438 2 134926 856
rect 135094 2 136582 856
rect 136750 2 138330 856
rect 138498 2 139986 856
rect 140154 2 141734 856
rect 141902 2 143390 856
rect 143558 2 145138 856
rect 145306 2 146794 856
rect 146962 2 148542 856
rect 148710 2 150198 856
rect 150366 2 151946 856
rect 152114 2 153602 856
rect 153770 2 155350 856
rect 155518 2 157006 856
rect 157174 2 158662 856
rect 158830 2 160410 856
rect 160578 2 162066 856
rect 162234 2 163814 856
rect 163982 2 165470 856
rect 165638 2 167218 856
rect 167386 2 168874 856
rect 169042 2 170622 856
rect 170790 2 172278 856
rect 172446 2 174026 856
rect 174194 2 175682 856
rect 175850 2 177430 856
rect 177598 2 179086 856
<< obsm3 >>
rect 841 35 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 62619 2048 65568 26485
rect 66048 2048 80928 26485
rect 81408 2048 96288 26485
rect 96768 2048 111648 26485
rect 112128 2048 121197 26485
rect 62619 443 121197 2048
<< labels >>
rlabel metal4 s 19568 2128 19888 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 VGND
port 1 nsew ground input
rlabel metal4 s 4208 2128 4528 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 VPWR
port 2 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 VPWR
port 2 nsew power input
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 4 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 5 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[0]
port 6 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[10]
port 7 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[11]
port 8 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[12]
port 9 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[13]
port 10 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[14]
port 11 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 wbs_adr_i[15]
port 12 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[16]
port 13 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[17]
port 14 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[18]
port 15 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_adr_i[19]
port 16 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[1]
port 17 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_adr_i[20]
port 18 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[21]
port 19 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 wbs_adr_i[22]
port 20 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 wbs_adr_i[23]
port 21 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 wbs_adr_i[24]
port 22 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_adr_i[25]
port 23 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 wbs_adr_i[26]
port 24 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 wbs_adr_i[27]
port 25 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 wbs_adr_i[28]
port 26 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 wbs_adr_i[29]
port 27 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[2]
port 28 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 wbs_adr_i[30]
port 29 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 wbs_adr_i[31]
port 30 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[3]
port 31 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[4]
port 32 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[5]
port 33 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[6]
port 34 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[7]
port 35 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[8]
port 36 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[9]
port 37 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_cyc_i
port 38 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[0]
port 39 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_i[10]
port 40 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_i[11]
port 41 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[12]
port 42 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_i[13]
port 43 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_i[14]
port 44 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[15]
port 45 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_dat_i[16]
port 46 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[17]
port 47 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wbs_dat_i[18]
port 48 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_i[19]
port 49 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[1]
port 50 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[20]
port 51 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[21]
port 52 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[22]
port 53 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_i[23]
port 54 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 wbs_dat_i[24]
port 55 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_i[25]
port 56 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 wbs_dat_i[26]
port 57 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 wbs_dat_i[27]
port 58 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 wbs_dat_i[28]
port 59 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 wbs_dat_i[29]
port 60 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[2]
port 61 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 wbs_dat_i[30]
port 62 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_i[31]
port 63 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[3]
port 64 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[4]
port 65 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[5]
port 66 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[6]
port 67 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[7]
port 68 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[8]
port 69 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[9]
port 70 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[0]
port 71 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[10]
port 72 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 wbs_dat_o[11]
port 73 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[12]
port 74 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[13]
port 75 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[14]
port 76 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_o[15]
port 77 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[16]
port 78 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_o[17]
port 79 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[18]
port 80 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_o[19]
port 81 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[1]
port 82 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 wbs_dat_o[20]
port 83 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 wbs_dat_o[21]
port 84 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 wbs_dat_o[22]
port 85 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_o[23]
port 86 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 wbs_dat_o[24]
port 87 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 wbs_dat_o[25]
port 88 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 wbs_dat_o[26]
port 89 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 wbs_dat_o[27]
port 90 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 wbs_dat_o[28]
port 91 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 wbs_dat_o[29]
port 92 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[2]
port 93 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 wbs_dat_o[30]
port 94 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 wbs_dat_o[31]
port 95 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[3]
port 96 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[4]
port 97 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[5]
port 98 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[6]
port 99 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[7]
port 100 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[8]
port 101 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[9]
port 102 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_sel_i[0]
port 103 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[1]
port 104 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_sel_i[2]
port 105 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_sel_i[3]
port 106 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_stb_i
port 107 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_we_i
port 108 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10654836
string GDS_FILE /mnt/c/Users/Ismael/Efabless-wsl/caravel_tutorial/caravel_example/openlane/SPM_example/runs/SPM_example/results/finishing/SPM_example.magic.gds
string GDS_START 476124
<< end >>

