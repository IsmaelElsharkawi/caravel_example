* NGSPICE file created from SPM_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt SPM_example VGND VPWR wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2106_ _2213_/A VGND VGND VPWR VPWR _2194_/A sky130_fd_sc_hd__buf_2
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2037_ _2285_/A VGND VGND VPWR VPWR _2083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2173__A2 _2118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1270_ _1268_/X _1263_/X _1269_/Y VGND VGND VPWR VPWR _1270_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1606_ _2445_/Q _2444_/Q _1606_/C VGND VGND VPWR VPWR _1612_/C sky130_fd_sc_hd__and3_1
X_2586_ _2595_/CLK _2586_/D _2350_/Y VGND VGND VPWR VPWR _2586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2164__A2 _2118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1537_ input48/X _2429_/Q _1545_/S VGND VGND VPWR VPWR _1538_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1468_ _1468_/A VGND VGND VPWR VPWR _2469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1399_ _1399_/A VGND VGND VPWR VPWR _2500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2185__A _2185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2522__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2440_ _2599_/CLK _2440_/D _1923_/Y VGND VGND VPWR VPWR _2440_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2371_ _2599_/CLK _2371_/D _1837_/Y VGND VGND VPWR VPWR _2371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1322_ _1320_/X _1313_/X _1321_/Y VGND VGND VPWR VPWR _1322_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1253_ input49/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1184_ _1184_/A _1184_/B VGND VGND VPWR VPWR _1187_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2545__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2137__A2 _2135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2569_ _2569_/CLK _2569_/D _2328_/Y VGND VGND VPWR VPWR _2569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1229__B1_N _1224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input55_A wbs_dat_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2418__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1940_ _1943_/A VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2272__B _2477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1871_ _1875_/A VGND VGND VPWR VPWR _1871_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2568__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1169__A _2013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2423_ _2576_/CLK _2423_/D _1902_/Y VGND VGND VPWR VPWR _2423_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2354_ _2354_/A VGND VGND VPWR VPWR _2354_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1305_ _1293_/X _1288_/X _1304_/Y VGND VGND VPWR VPWR _1305_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2285_ _2285_/A _2285_/B _2438_/Q VGND VGND VPWR VPWR _2285_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1236_ _2247_/A VGND VGND VPWR VPWR _2024_/B sky130_fd_sc_hd__buf_2
XFILLER_42_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1167_ _1167_/A _1167_/B VGND VGND VPWR VPWR _1168_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _2519_/Q VGND VGND VPWR VPWR _2070_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _1925_/A VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1854_ _1856_/A VGND VGND VPWR VPWR _1854_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1548__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1785_ _2589_/Q _2586_/Q _1784_/B VGND VGND VPWR VPWR _2589_/D sky130_fd_sc_hd__a21o_1
XFILLER_11_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2406_ _2549_/CLK _2406_/D _1880_/Y VGND VGND VPWR VPWR _2406_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2337_ _2355_/A VGND VGND VPWR VPWR _2342_/A sky130_fd_sc_hd__buf_2
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2268_ _2264_/Y _2266_/Y _2267_/X VGND VGND VPWR VPWR _2268_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1219_ _1297_/A VGND VGND VPWR VPWR _1219_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1512__D _1512_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2199_ _2500_/Q _2198_/X _2165_/X _2189_/X VGND VGND VPWR VPWR _2199_/X sky130_fd_sc_hd__o31a_1
XFILLER_22_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1272__A _1297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input18_A wbs_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1570_ input63/X _2414_/Q _1578_/S VGND VGND VPWR VPWR _1571_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2278__A _2285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1182__A _1182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2165_/A VGND VGND VPWR VPWR _2122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2053_ _2083_/A _2061_/B _2411_/Q VGND VGND VPWR VPWR _2053_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_48_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1910__A _1912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1906_ _1906_/A VGND VGND VPWR VPWR _1906_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1837_ _1838_/A VGND VGND VPWR VPWR _1837_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1768_ _2585_/Q _2582_/Q VGND VGND VPWR VPWR _1768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1699_ _1696_/X _1697_/Y _1706_/C _2414_/Q VGND VGND VPWR VPWR _1700_/B sky130_fd_sc_hd__and4bb_1
XFILLER_85_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 _2528_/Q VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput86 _2538_/Q VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput97 _2519_/Q VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _1622_/A _1622_/B VGND VGND VPWR VPWR _2370_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1553_ _1553_/A VGND VGND VPWR VPWR _2422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1484_ _2461_/Q _2462_/Q _1484_/S VGND VGND VPWR VPWR _1485_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2105_ _2523_/Q VGND VGND VPWR VPWR _2105_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2036_ _2515_/Q VGND VGND VPWR VPWR _2036_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2100__B1 _2074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2451__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2291__A _2545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1605_ _1586_/B _1606_/C _1604_/Y VGND VGND VPWR VPWR _2444_/D sky130_fd_sc_hd__a21oi_1
XFILLER_173_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2585_ _2595_/CLK _2585_/D _2348_/Y VGND VGND VPWR VPWR _2585_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1536_ _1558_/A VGND VGND VPWR VPWR _1545_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1467_ _2469_/Q _2470_/Q _1473_/S VGND VGND VPWR VPWR _1468_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1398_ _2500_/Q _2501_/Q _1406_/S VGND VGND VPWR VPWR _1399_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2474__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2185__B _2228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2019_ _2026_/A _2252_/A VGND VGND VPWR VPWR _2231_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2370_ _2599_/CLK _2370_/D _1836_/Y VGND VGND VPWR VPWR _2370_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1321_ _2555_/Q VGND VGND VPWR VPWR _1321_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1252_ _1374_/A VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2497__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2286__A _2294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1183_ _1183_/A input9/X VGND VGND VPWR VPWR _1187_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1621__C _1621_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1365__A _2546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2568_ _2576_/CLK _2568_/D _2327_/Y VGND VGND VPWR VPWR _2568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1345__A1 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1519_ input56/X _2437_/Q _1523_/S VGND VGND VPWR VPWR _1520_/A sky130_fd_sc_hd__mux2_1
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2499_ _2512_/CLK _2499_/D _1996_/Y VGND VGND VPWR VPWR _2499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2196__A _2229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input48_A wbs_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1870_ _1882_/A VGND VGND VPWR VPWR _1875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2422_ _2512_/CLK _2422_/D _1900_/Y VGND VGND VPWR VPWR _2422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2353_ _2354_/A VGND VGND VPWR VPWR _2353_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1913__A _1913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1304_ _2558_/Q VGND VGND VPWR VPWR _1304_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2284_ _2544_/Q VGND VGND VPWR VPWR _2284_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1235_ _2026_/A VGND VGND VPWR VPWR _2247_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1166_ _1166_/A _1166_/B VGND VGND VPWR VPWR _1168_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2055__A2 _2292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2512__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1999_ _1999_/A VGND VGND VPWR VPWR _1999_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2535__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _1925_/A VGND VGND VPWR VPWR _1922_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1853_ _1856_/A VGND VGND VPWR VPWR _1853_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1908__A _1912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1784_ _1784_/A _1784_/B VGND VGND VPWR VPWR _2588_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2405_ _2595_/CLK _2405_/D _1879_/Y VGND VGND VPWR VPWR _2405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1643__A _1643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2336_ _2336_/A VGND VGND VPWR VPWR _2336_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2267_ _2508_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2267_/X sky130_fd_sc_hd__o31a_1
XFILLER_6_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1218_ _2237_/A VGND VGND VPWR VPWR _1297_/A sky130_fd_sc_hd__buf_2
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2276__A2 _2246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2198_ _2241_/A VGND VGND VPWR VPWR _2198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2408__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2558__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2278__B _2285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2121_ _1673_/C _2118_/X _2119_/X _2120_/Y VGND VGND VPWR VPWR _2121_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2052_ _2517_/Q VGND VGND VPWR VPWR _2052_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2294__A _2294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1905_ _1906_/A VGND VGND VPWR VPWR _1905_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1836_ _1838_/A VGND VGND VPWR VPWR _1836_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1767_ _2585_/Q _2582_/Q VGND VGND VPWR VPWR _1767_/X sky130_fd_sc_hd__and2_1
XFILLER_190_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1698_ _1647_/X _2414_/Q _1696_/X _1697_/Y VGND VGND VPWR VPWR _1700_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2319_ _2323_/A VGND VGND VPWR VPWR _2319_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2380__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput76 _2529_/Q VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 _2539_/Q VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_81_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput98 _2520_/Q VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2098__B _2161_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_A wbs_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2024__C_N _2408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1621_ _1643_/A _1621_/B _1621_/C _1621_/D VGND VGND VPWR VPWR _1622_/B sky130_fd_sc_hd__nor4_1
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1552_ input40/X _2422_/Q _1556_/S VGND VGND VPWR VPWR _1553_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1483_ _1483_/A VGND VGND VPWR VPWR _2462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1193__A _2448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2104_ _2097_/Y _2071_/X _2103_/Y VGND VGND VPWR VPWR _2522_/D sky130_fd_sc_hd__o21ai_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2035_ _2018_/Y _2022_/X _2034_/Y VGND VGND VPWR VPWR _2514_/D sky130_fd_sc_hd__o21ai_2
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2100__A1 _1686_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1819_ _2601_/Q _2598_/Q VGND VGND VPWR VPWR _1819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2167__A1 _2161_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1831__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1604_ _1586_/B _1606_/C _1194_/X VGND VGND VPWR VPWR _1604_/Y sky130_fd_sc_hd__o21ai_1
X_2584_ _2595_/CLK _2584_/D _2347_/Y VGND VGND VPWR VPWR _2584_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1535_ _1535_/A VGND VGND VPWR VPWR _2430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1466_ _1466_/A VGND VGND VPWR VPWR _2470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1397_ _1430_/A VGND VGND VPWR VPWR _1406_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1651__A _2546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2018_ _2514_/Q VGND VGND VPWR VPWR _2018_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2085__B1 _2074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1363__A2 _1339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2076__B1 _2074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1500__S _1506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1736__A _2546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1354__A2 _1339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1320_ _1346_/A VGND VGND VPWR VPWR _1320_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1251_ _1497_/A VGND VGND VPWR VPWR _1374_/A sky130_fd_sc_hd__buf_2
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1182_ _1182_/A _1182_/B _1182_/C VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1801__A1_N _1652_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_wb_clk_i clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1646__A _2546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2567_ _2576_/CLK _2567_/D _2326_/Y VGND VGND VPWR VPWR _2567_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1518_ _1518_/A VGND VGND VPWR VPWR _2438_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2441__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2498_ _2512_/CLK _2498_/D _1995_/Y VGND VGND VPWR VPWR _2498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1449_ _2477_/Q _2478_/Q _1451_/S VGND VGND VPWR VPWR _1450_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2591__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2230__B1 _2205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2049__B1 _2246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2464__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2421_ _2512_/CLK _2421_/D _1899_/Y VGND VGND VPWR VPWR _2421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2352_ _2354_/A VGND VGND VPWR VPWR _2352_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1303_ input38/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1303_/X sky130_fd_sc_hd__o21ba_1
X_2283_ _2277_/Y _2246_/X _2282_/Y VGND VGND VPWR VPWR _2543_/D sky130_fd_sc_hd__o21ai_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1234_ input52/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1234_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2288__B1 _2032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1165_ _1165_/A _1165_/B VGND VGND VPWR VPWR _1165_/Y sky130_fd_sc_hd__nand2_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1998_ _1999_/A VGND VGND VPWR VPWR _1998_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2000__A _2006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2487__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1286__A _1608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input60_A wbs_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1921_ _1925_/A VGND VGND VPWR VPWR _1921_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1852_ _1856_/A VGND VGND VPWR VPWR _1852_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1783_ _1780_/X _1781_/Y _1789_/C _2433_/Q VGND VGND VPWR VPWR _1784_/B sky130_fd_sc_hd__and4bb_1
XFILLER_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2404_ _2595_/CLK _2404_/D _1878_/Y VGND VGND VPWR VPWR _2404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2335_ _2336_/A VGND VGND VPWR VPWR _2335_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2266_ _1226_/Y _2237_/X _2249_/X _2265_/Y VGND VGND VPWR VPWR _2266_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_6_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1217_ _2576_/Q _1209_/X _1211_/X _1216_/Y VGND VGND VPWR VPWR _2575_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2197_ _1269_/Y _2135_/X _2162_/X _2196_/Y VGND VGND VPWR VPWR _2197_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_26_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2502__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2120_ _2144_/A _2459_/Q VGND VGND VPWR VPWR _2120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2051_ _2045_/Y _2022_/X _2050_/Y VGND VGND VPWR VPWR _2516_/D sky130_fd_sc_hd__o21ai_1
XFILLER_130_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1919__A _2361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1904_ _1906_/A VGND VGND VPWR VPWR _1904_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1835_ _1838_/A VGND VGND VPWR VPWR _1835_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1766_ _2583_/Q _2580_/Q _1765_/B VGND VGND VPWR VPWR _2583_/D sky130_fd_sc_hd__a21o_1
XFILLER_50_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1697_ _2393_/Q _2390_/Q VGND VGND VPWR VPWR _1697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2324_/A VGND VGND VPWR VPWR _2323_/A sky130_fd_sc_hd__buf_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2249_ _2249_/A VGND VGND VPWR VPWR _2249_/X sky130_fd_sc_hd__buf_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2525__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput77 _2530_/Q VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput88 _2540_/Q VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 _2521_/Q VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_172_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input23_A wbs_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1620_ _1828_/A _1621_/C _1621_/D _1621_/B VGND VGND VPWR VPWR _1622_/A sky130_fd_sc_hd__o22a_1
XANTENNA_output91_A _2543_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1551_ _1551_/A VGND VGND VPWR VPWR _2423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1482_ _2462_/Q _2463_/Q _1484_/S VGND VGND VPWR VPWR _1483_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2103_ _2098_/Y _2100_/Y _2102_/X VGND VGND VPWR VPWR _2103_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2034_ _2024_/Y _2031_/Y _2033_/Y VGND VGND VPWR VPWR _2034_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2100__A2 _1583_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2548__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1818_ _2601_/Q _2598_/Q VGND VGND VPWR VPWR _1818_/X sky130_fd_sc_hd__and2_1
XFILLER_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1749_ _2579_/Q _2404_/Q VGND VGND VPWR VPWR _1749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1815__C _1815_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2562__RESET_B _2320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1188__B _1188_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1603_ _1603_/A VGND VGND VPWR VPWR _2443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2583_ _2595_/CLK _2583_/D _2346_/Y VGND VGND VPWR VPWR _2583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1534_ input49/X _2430_/Q _1534_/S VGND VGND VPWR VPWR _1535_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1465_ _2470_/Q _2471_/Q _1473_/S VGND VGND VPWR VPWR _1466_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ _1396_/A VGND VGND VPWR VPWR _2501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2017_ _1214_/X _2016_/X _2513_/Q VGND VGND VPWR VPWR _2513_/D sky130_fd_sc_hd__a21oi_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2370__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2003__A _2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ _2570_/Q _1233_/X _1247_/X _1249_/Y VGND VGND VPWR VPWR _2569_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1181_ input4/X input3/X VGND VGND VPWR VPWR _1182_/C sky130_fd_sc_hd__nor2_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1814__A1 _1722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1578__A0 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2566_ _2576_/CLK _2566_/D _2325_/Y VGND VGND VPWR VPWR _2566_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1517_ input58/X _2438_/Q _1523_/S VGND VGND VPWR VPWR _1518_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2497_ _2512_/CLK _2497_/D _1993_/Y VGND VGND VPWR VPWR _2497_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1448_ _1448_/A VGND VGND VPWR VPWR _2478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1379_ _2508_/Q _2509_/Q _1383_/S VGND VGND VPWR VPWR _1380_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1747__A _1747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2420_ _2560_/CLK _2420_/D _1898_/Y VGND VGND VPWR VPWR _2420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2351_ _2354_/A VGND VGND VPWR VPWR _2351_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1302_ _1374_/A VGND VGND VPWR VPWR _1302_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2282_ _2278_/Y _2280_/Y _2281_/X VGND VGND VPWR VPWR _2282_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ _1608_/B VGND VGND VPWR VPWR _1233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1164_ _1200_/A VGND VGND VPWR VPWR _2213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ _1999_/A VGND VGND VPWR VPWR _1997_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2549_ _2549_/CLK _2549_/D _2304_/Y VGND VGND VPWR VPWR _2549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input53_A wbs_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1506__S _1506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1733__C _1751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ _1944_/A VGND VGND VPWR VPWR _1925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_143_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2431__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ _2367_/A VGND VGND VPWR VPWR _1856_/A sky130_fd_sc_hd__buf_2
XFILLER_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1782_ _1747_/X _2433_/Q _1780_/X _1781_/Y VGND VGND VPWR VPWR _1784_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2581__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2403_ _2459_/CLK _2403_/D _1877_/Y VGND VGND VPWR VPWR _2403_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2334_ _2336_/A VGND VGND VPWR VPWR _2334_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2265_ _2272_/A _2476_/Q VGND VGND VPWR VPWR _2265_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1216_ _1212_/X _1214_/X _1215_/Y VGND VGND VPWR VPWR _1216_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2196_ _2229_/A _2468_/Q VGND VGND VPWR VPWR _2196_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2011__A _2011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2454__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1227__A2 _1214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1297__A _1297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2050_ _2046_/Y _2048_/Y _2049_/X VGND VGND VPWR VPWR _2050_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_130_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1903_ _1906_/A VGND VGND VPWR VPWR _1903_/Y sky130_fd_sc_hd__inv_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ _1838_/A VGND VGND VPWR VPWR _1834_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1765_ _1765_/A _1765_/B VGND VGND VPWR VPWR _2582_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1696_ _2393_/Q _2390_/Q VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__and2_1
XFILLER_172_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2317_/A VGND VGND VPWR VPWR _2317_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2477__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2264_/A _2285_/B _2433_/Q VGND VGND VPWR VPWR _2248_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2179_ _2187_/A _2466_/Q VGND VGND VPWR VPWR _2179_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2006__A _2006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 _2531_/Q VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 _2541_/Q VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1580__A _2186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A wbs_adr_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1620__A2 _1621_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ input41/X _2423_/Q _1556_/S VGND VGND VPWR VPWR _1551_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1481_ _1481_/A VGND VGND VPWR VPWR _2463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2102_ _2489_/Q _2066_/X _2078_/X _2101_/X VGND VGND VPWR VPWR _2102_/X sky130_fd_sc_hd__o31a_1
XFILLER_95_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2033_ _2481_/Q _2074_/A _2032_/X VGND VGND VPWR VPWR _2033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1817_ _2599_/Q _2596_/Q _1816_/B VGND VGND VPWR VPWR _2599_/D sky130_fd_sc_hd__a21o_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1748_ _2579_/Q _2404_/Q VGND VGND VPWR VPWR _1748_/X sky130_fd_sc_hd__and2_1
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1679_ _1676_/X _1677_/Y _1706_/C _2417_/Q VGND VGND VPWR VPWR _1680_/B sky130_fd_sc_hd__and4bb_1
XFILLER_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input8_A wbs_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2094__A2 _2066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1602_ _1606_/C _1614_/C _1602_/C VGND VGND VPWR VPWR _1603_/A sky130_fd_sc_hd__and3b_1
X_2582_ _2595_/CLK _2582_/D _2345_/Y VGND VGND VPWR VPWR _2582_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1533_ _1533_/A VGND VGND VPWR VPWR _2431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1464_ _1486_/A VGND VGND VPWR VPWR _1473_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ _2501_/Q _2502_/Q _1395_/S VGND VGND VPWR VPWR _1396_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2016_ _2252_/A VGND VGND VPWR VPWR _2016_/X sky130_fd_sc_hd__buf_2
XFILLER_24_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2085__A2 _2062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2515__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1211__B1_N _1339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2076__A2 _2062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1284__B1 _2171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1182_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2538__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2067__A2 _2066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1275__B1 _2185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1814__A2 _1815_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2565_ _2576_/CLK _2565_/D _2323_/Y VGND VGND VPWR VPWR _2565_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1516_ _1516_/A VGND VGND VPWR VPWR _2439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2496_ _2512_/CLK _2496_/D _1992_/Y VGND VGND VPWR VPWR _2496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1447_ _2478_/Q _2479_/Q _1451_/S VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1378_ _1378_/A VGND VGND VPWR VPWR _2509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2230__A2 _2186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2014__A _2014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2350_ _2354_/A VGND VGND VPWR VPWR _2350_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1301_ _2560_/Q _1286_/X _1298_/X _1300_/Y VGND VGND VPWR VPWR _2559_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2281_ _2510_/Q _2066_/A _2252_/X _2032_/X VGND VGND VPWR VPWR _2281_/X sky130_fd_sc_hd__o31a_1
XFILLER_26_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1232_ _2573_/Q _1209_/X _1229_/X _1231_/Y VGND VGND VPWR VPWR _2572_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2288__A2 _2066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _1999_/A VGND VGND VPWR VPWR _1996_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1673__A _1777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2548_ _2553_/CLK _2548_/D _2303_/Y VGND VGND VPWR VPWR _2548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2479_ _2512_/CLK _2479_/D _1971_/Y VGND VGND VPWR VPWR _2479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2009__A _2011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2383__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A wbs_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1733__D _2409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1850_ _1850_/A VGND VGND VPWR VPWR _1850_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1781_ _2589_/Q _2586_/Q VGND VGND VPWR VPWR _1781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2402_ _2459_/CLK _2402_/D _1875_/Y VGND VGND VPWR VPWR _2402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2333_ _2336_/A VGND VGND VPWR VPWR _2333_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2264_ _2264_/A _2285_/B _2435_/Q VGND VGND VPWR VPWR _2264_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1215_ _2575_/Q VGND VGND VPWR VPWR _1215_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2195_ _2238_/A VGND VGND VPWR VPWR _2229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1979_ _1980_/A VGND VGND VPWR VPWR _1979_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2121__A1 _1673_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2188__A1 _1828_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1744__C _1751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1902_ _1906_/A VGND VGND VPWR VPWR _1902_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1833_ _2367_/A VGND VGND VPWR VPWR _1838_/A sky130_fd_sc_hd__buf_2
XFILLER_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1764_ _1761_/X _1762_/Y _1789_/C _2436_/Q VGND VGND VPWR VPWR _1765_/B sky130_fd_sc_hd__and4bb_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1695_ _2391_/Q _2388_/Q _1694_/B VGND VGND VPWR VPWR _2391_/D sky130_fd_sc_hd__a21o_1
XFILLER_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1951__A _1975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2317_/A VGND VGND VPWR VPWR _2316_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2247_ _2247_/A VGND VGND VPWR VPWR _2285_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ _2178_/A _2228_/B VGND VGND VPWR VPWR _2178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2022__A _2116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput79 _2532_/Q VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2421__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2571__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1480_ _2463_/Q _2464_/Q _1484_/S VGND VGND VPWR VPWR _1481_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2101_ _2146_/A VGND VGND VPWR VPWR _2101_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2032_ _2231_/A VGND VGND VPWR VPWR _2032_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2107__A _2194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1816_ _1816_/A _1816_/B VGND VGND VPWR VPWR _2598_/D sky130_fd_sc_hd__nor2_1
XFILLER_15_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1747_ _1747_/A VGND VGND VPWR VPWR _1747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2444__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1678_ _1647_/X _2417_/Q _1676_/X _1677_/Y VGND VGND VPWR VPWR _1680_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2594__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2094__A3 _2078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2467__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1601_ _1588_/A _1593_/A _2442_/Q _2443_/Q VGND VGND VPWR VPWR _1602_/C sky130_fd_sc_hd__a31o_1
XFILLER_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2581_ _2595_/CLK _2581_/D _2344_/Y VGND VGND VPWR VPWR _2581_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1532_ input50/X _2431_/Q _1534_/S VGND VGND VPWR VPWR _1533_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1463_ _1463_/A VGND VGND VPWR VPWR _2471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1394_ _1394_/A VGND VGND VPWR VPWR _2502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2015_ _2028_/B _2028_/C _2028_/D VGND VGND VPWR VPWR _2252_/A sky130_fd_sc_hd__nand3_4
XFILLER_110_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2300__A _2324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2067__A3 _2016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2564_ _2576_/CLK _2564_/D _2322_/Y VGND VGND VPWR VPWR _2564_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1515_ input59/X _2439_/Q _1523_/S VGND VGND VPWR VPWR _1516_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2495_ _2512_/CLK _2495_/D _1991_/Y VGND VGND VPWR VPWR _2495_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1435__S _1439_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2120__A _2144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1446_ _1446_/A VGND VGND VPWR VPWR _2479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1377_ _2509_/Q _2510_/Q _1383_/S VGND VGND VPWR VPWR _1378_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2030__A _2074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2049__A3 _2016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1257__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2205__A _2249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2505__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1300_ _1293_/X _1288_/X _1299_/Y VGND VGND VPWR VPWR _1300_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2280_ _1215_/Y _2237_/X _2249_/X _2279_/Y VGND VGND VPWR VPWR _2280_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1231_ _1212_/X _1214_/X _2257_/A VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1995_ _1999_/A VGND VGND VPWR VPWR _1995_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1225__B1_N _1224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2547_ _2549_/CLK _2547_/D _2302_/Y VGND VGND VPWR VPWR _2547_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2478_ _2512_/CLK _2478_/D _1970_/Y VGND VGND VPWR VPWR _2478_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1429_ _1429_/A VGND VGND VPWR VPWR _2486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2025__A _2237_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2528__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A wbs_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1780_ _2589_/Q _2586_/Q VGND VGND VPWR VPWR _1780_/X sky130_fd_sc_hd__and2_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2401_ _2459_/CLK _2401_/D _1874_/Y VGND VGND VPWR VPWR _2401_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2332_ _2336_/A VGND VGND VPWR VPWR _2332_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2263_ _2541_/Q VGND VGND VPWR VPWR _2263_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1214_ _2054_/A VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__buf_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2194_ _2194_/A _2236_/B _2427_/Q VGND VGND VPWR VPWR _2194_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_22_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ _1980_/A VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2197__A2 _2135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2271__C_N _2436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2599_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2121__A2 _2118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2188__A2 _2186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1744__D _2408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _1913_/A VGND VGND VPWR VPWR _1906_/A sky130_fd_sc_hd__buf_2
XFILLER_203_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1832_ _2361_/A VGND VGND VPWR VPWR _2367_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1763_ _1747_/X _2436_/Q _1761_/X _1762_/Y VGND VGND VPWR VPWR _1765_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_184_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1694_ _1694_/A _1694_/B VGND VGND VPWR VPWR _2390_/D sky130_fd_sc_hd__nor2_1
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2317_/A VGND VGND VPWR VPWR _2315_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2246_/A VGND VGND VPWR VPWR _2246_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2177_ _2531_/Q VGND VGND VPWR VPWR _2177_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2373__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2303__A _2305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput69 _2513_/Q VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_81_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1550__A0 input41/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1589__A _1589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2213__A _2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2100_ _1686_/C _1583_/S _2074_/X _2099_/Y VGND VGND VPWR VPWR _2100_/Y sky130_fd_sc_hd__o211ai_1
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2031_ _1672_/A _2292_/B _2027_/Y _2030_/X VGND VGND VPWR VPWR _2031_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2107__B _2134_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1815_ _1828_/A _1815_/B _1815_/C _1815_/D VGND VGND VPWR VPWR _1816_/B sky130_fd_sc_hd__nor4_1
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1746_ _2407_/Q _2402_/Q _1745_/B VGND VGND VPWR VPWR _2407_/D sky130_fd_sc_hd__a21o_1
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1677_ _2387_/Q _2384_/Q VGND VGND VPWR VPWR _1677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1532__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2229_ _2229_/A _2472_/Q VGND VGND VPWR VPWR _2229_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1202__A _2241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1523__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A wbs_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2208__A _2252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ _2441_/Q _2440_/Q _2443_/Q _2442_/Q VGND VGND VPWR VPWR _1606_/C sky130_fd_sc_hd__and4_1
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2580_ _2595_/CLK _2580_/D _2342_/Y VGND VGND VPWR VPWR _2580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1531_ _1531_/A VGND VGND VPWR VPWR _2432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1462_ _2471_/Q _2472_/Q _1462_/S VGND VGND VPWR VPWR _1463_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1393_ _2502_/Q _2503_/Q _1395_/S VGND VGND VPWR VPWR _1394_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2014_ _2014_/A _2014_/B VGND VGND VPWR VPWR _2028_/D sky130_fd_sc_hd__nor2_4
XFILLER_3_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2118__A _2186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1957__A _1975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2411__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1729_ _2401_/Q _2398_/Q _1728_/B VGND VGND VPWR VPWR _2401_/D sky130_fd_sc_hd__a21o_1
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2561__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2028__A _2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1777__A _1777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2584__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2563_ _2576_/CLK _2563_/D _2321_/Y VGND VGND VPWR VPWR _2563_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1514_ _1558_/A VGND VGND VPWR VPWR _1523_/S sky130_fd_sc_hd__buf_2
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2494_ _2512_/CLK _2494_/D _1990_/Y VGND VGND VPWR VPWR _2494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1445_ _2479_/Q _2480_/Q _1451_/S VGND VGND VPWR VPWR _1446_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1376_ _1376_/A VGND VGND VPWR VPWR _2510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2221__A _2264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _2572_/Q VGND VGND VPWR VPWR _2257_/A sky130_fd_sc_hd__inv_2
XFILLER_133_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1994_ _2006_/A VGND VGND VPWR VPWR _1999_/A sky130_fd_sc_hd__buf_2
XFILLER_33_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1673__C _1673_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2546_ _2549_/CLK _2546_/D _2301_/Y VGND VGND VPWR VPWR _2546_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2477_ _2595_/CLK _2477_/D _1968_/Y VGND VGND VPWR VPWR _2477_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1428_ _2486_/Q _2487_/Q _1428_/S VGND VGND VPWR VPWR _1429_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1359_ _2549_/Q _1339_/X _1356_/X _1358_/Y VGND VGND VPWR VPWR _2548_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2306__A _2324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1880__A _1881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ _2459_/CLK _2400_/D _1873_/Y VGND VGND VPWR VPWR _2400_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2331_ _2355_/A VGND VGND VPWR VPWR _2336_/A sky130_fd_sc_hd__buf_2
XFILLER_152_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2262_ _2256_/Y _2246_/X _2261_/Y VGND VGND VPWR VPWR _2540_/D sky130_fd_sc_hd__o21ai_1
XFILLER_152_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1213_ _2238_/A VGND VGND VPWR VPWR _2054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2193_ _2533_/Q VGND VGND VPWR VPWR _2193_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1977_ _1980_/A VGND VGND VPWR VPWR _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2529_ _2569_/CLK _2529_/D VGND VGND VPWR VPWR _2529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1205__A _2238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2036__A _2515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input51_A wbs_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2112__A3 _2078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ _1900_/A VGND VGND VPWR VPWR _1900_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1831_ input1/X VGND VGND VPWR VPWR _2361_/A sky130_fd_sc_hd__buf_2
XFILLER_54_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1762_ _2583_/Q _2580_/Q VGND VGND VPWR VPWR _1762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1693_ _1777_/A _1693_/B _1693_/C _1693_/D VGND VGND VPWR VPWR _1694_/B sky130_fd_sc_hd__nor4_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2314_ _2317_/A VGND VGND VPWR VPWR _2314_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _2539_/Q VGND VGND VPWR VPWR _2245_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2176_ _2169_/Y _2160_/X _2175_/Y VGND VGND VPWR VPWR _2530_/D sky130_fd_sc_hd__o21ai_1
XFILLER_211_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2518__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2030_ _2074_/A VGND VGND VPWR VPWR _2030_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1814_ _1722_/X _1815_/C _1815_/D _1815_/B VGND VGND VPWR VPWR _1816_/A sky130_fd_sc_hd__o22a_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1745_ _1745_/A _1745_/B VGND VGND VPWR VPWR _2406_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _2387_/Q _2384_/Q VGND VGND VPWR VPWR _1676_/X sky130_fd_sc_hd__and2_1
XFILLER_171_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2228_ _2228_/A _2228_/B VGND VGND VPWR VPWR _2228_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2088__A2 _2071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _2529_/Q VGND VGND VPWR VPWR _2159_/Y sky130_fd_sc_hd__inv_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2490__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2314__A _2317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1523__A1 _2435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2079__A2 _2066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wbs_adr_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1530_ input51/X _2432_/Q _1534_/S VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1461_ _1461_/A VGND VGND VPWR VPWR _2472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1392_ _1392_/A VGND VGND VPWR VPWR _2503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2013_ _2013_/A _2013_/B VGND VGND VPWR VPWR _2014_/B sky130_fd_sc_hd__nand2_2
XFILLER_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2134__A _2194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1728_ _1728_/A _1728_/B VGND VGND VPWR VPWR _2400_/D sky130_fd_sc_hd__nor2_1
XFILLER_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1168__A_N _1165_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1659_ _1655_/X _1656_/Y _1706_/C _2420_/Q VGND VGND VPWR VPWR _1660_/B sky130_fd_sc_hd__and4bb_1
XFILLER_63_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input6_A wbs_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1213__A _2238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2028__B _2028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2386__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2562_ _2576_/CLK _2562_/D _2320_/Y VGND VGND VPWR VPWR _2562_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1513_ _2186_/A VGND VGND VPWR VPWR _1558_/A sky130_fd_sc_hd__buf_2
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2493_ _2512_/CLK _2493_/D _1989_/Y VGND VGND VPWR VPWR _2493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1444_ _1444_/A VGND VGND VPWR VPWR _2480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1375_ _2510_/Q _2511_/Q _1383_/S VGND VGND VPWR VPWR _1376_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1726__A1 _1722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1208__A _1497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2039__A _2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1878__A _1881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2221__B _2236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2551__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1993_ _1993_/A VGND VGND VPWR VPWR _1993_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2545_ _2569_/CLK _2545_/D VGND VGND VPWR VPWR _2545_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_170_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2476_ _2512_/CLK _2476_/D _1967_/Y VGND VGND VPWR VPWR _2476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1427_ _1427_/A VGND VGND VPWR VPWR _2487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ _1346_/X _1341_/X _2046_/A VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1289_ _2561_/Q VGND VGND VPWR VPWR _2161_/A sky130_fd_sc_hd__inv_2
XFILLER_23_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2322__A _2323_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2424__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1372__S _1372_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2574__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1758__D _2437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2330_ input1/X VGND VGND VPWR VPWR _2355_/A sky130_fd_sc_hd__buf_2
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2261_ _2257_/Y _2259_/Y _2260_/X VGND VGND VPWR VPWR _2261_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1212_ _1293_/A VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2192_ _2184_/Y _2160_/X _2191_/Y VGND VGND VPWR VPWR _2532_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1311__A _1339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1976_ _1980_/A VGND VGND VPWR VPWR _1976_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2142__A _2247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2447__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1981__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2528_ _2560_/CLK _2528_/D VGND VGND VPWR VPWR _2528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2597__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2459_ _2459_/CLK _2459_/D _1946_/Y VGND VGND VPWR VPWR _2459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2317__A _2317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2042__B1 _2246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1891__A _1894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_A wbs_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2281__B1 _2032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ _2369_/Q _2600_/Q _1829_/B VGND VGND VPWR VPWR _2369_/D sky130_fd_sc_hd__a21o_1
XFILLER_19_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2033__B1 _2032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1761_ _2583_/Q _2580_/Q VGND VGND VPWR VPWR _1761_/X sky130_fd_sc_hd__and2_1
XFILLER_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1692_ _1631_/X _1693_/C _1693_/D _1693_/B VGND VGND VPWR VPWR _1694_/A sky130_fd_sc_hd__o22a_1
XFILLER_176_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2317_/A VGND VGND VPWR VPWR _2313_/Y sky130_fd_sc_hd__inv_2
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2235_/Y _2203_/X _2243_/Y VGND VGND VPWR VPWR _2538_/D sky130_fd_sc_hd__o21ai_1
XFILLER_41_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2549_/CLK sky130_fd_sc_hd__clkbuf_16
X_2175_ _2171_/Y _2173_/Y _2174_/X VGND VGND VPWR VPWR _2175_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1976__A _1980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1959_ _1962_/A VGND VGND VPWR VPWR _1959_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2047__A _2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1369__A2 _1194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1813_ _2599_/Q _2596_/Q VGND VGND VPWR VPWR _1815_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1744_ _1741_/X _1742_/Y _1751_/C _2408_/Q VGND VGND VPWR VPWR _1745_/B sky130_fd_sc_hd__and4bb_1
XFILLER_69_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1675_ _2385_/Q _2382_/Q _1674_/B VGND VGND VPWR VPWR _2385_/D sky130_fd_sc_hd__a21o_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2227_ _2537_/Q VGND VGND VPWR VPWR _2227_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _2150_/Y _2116_/X _2157_/Y VGND VGND VPWR VPWR _2528_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2089_ _2521_/Q VGND VGND VPWR VPWR _2089_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1220__A1 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2330__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2079__A3 _2078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1287__A1 input41/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1211__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2508__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1460_ _2472_/Q _2473_/Q _1462_/S VGND VGND VPWR VPWR _1461_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output75_A _2528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1391_ _2503_/Q _2504_/Q _1395_/S VGND VGND VPWR VPWR _1392_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2012_ _2448_/Q _2012_/B VGND VGND VPWR VPWR _2013_/B sky130_fd_sc_hd__nor2_1
XFILLER_188_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_32_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2134__B _2134_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1727_ _1777_/A _1727_/B _1727_/C _1727_/D VGND VGND VPWR VPWR _1728_/B sky130_fd_sc_hd__nor4_1
XFILLER_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2150__A _2528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1658_ _1747_/A VGND VGND VPWR VPWR _1706_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1589_ _1589_/A VGND VGND VPWR VPWR _1614_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2325__A _2329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1777__C _1777_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2561_ _2576_/CLK _2561_/D _2319_/Y VGND VGND VPWR VPWR _2561_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1512_ _1512_/A _2028_/B _2028_/C _1512_/D VGND VGND VPWR VPWR _2186_/A sky130_fd_sc_hd__nand4_4
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2492_ _2512_/CLK _2492_/D _1987_/Y VGND VGND VPWR VPWR _2492_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2480__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1443_ _2480_/Q _2481_/Q _1451_/S VGND VGND VPWR VPWR _1444_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1374_ _1374_/A VGND VGND VPWR VPWR _1383_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1984__A _1987_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1726__A2 _1727_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2559__RESET_B _2316_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1224__A _1589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2039__B _2450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1894__A _1894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1992_ _1993_/A VGND VGND VPWR VPWR _1992_/Y sky130_fd_sc_hd__inv_2
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2544_ _2569_/CLK _2544_/D VGND VGND VPWR VPWR _2544_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_118_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2475_ _2595_/CLK _2475_/D _1966_/Y VGND VGND VPWR VPWR _2475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1426_ _2487_/Q _2488_/Q _1428_/S VGND VGND VPWR VPWR _1427_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1357_ _2548_/Q VGND VGND VPWR VPWR _2046_/A sky130_fd_sc_hd__inv_2
XFILLER_25_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1288_ _2024_/B VGND VGND VPWR VPWR _1288_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1979__A _1980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2376__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1219__A _1297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1889__A _1913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1563__S _1567_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2260_ _2507_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2260_/X sky130_fd_sc_hd__o31a_1
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1211_ input56/X _1191_/X _1339_/A VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__o21ba_1
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2191_ _2185_/Y _2188_/Y _2190_/X VGND VGND VPWR VPWR _2191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1975_ _1975_/A VGND VGND VPWR VPWR _1980_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2527_ _2560_/CLK _2527_/D VGND VGND VPWR VPWR _2527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2458_ _2459_/CLK _2458_/D _1945_/Y VGND VGND VPWR VPWR _2458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1409_ _2495_/Q _2496_/Q _1417_/S VGND VGND VPWR VPWR _1410_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2389_ _2459_/CLK _2389_/D _1860_/Y VGND VGND VPWR VPWR _2389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2541__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input37_A wbs_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1760_ _2581_/Q _2578_/Q _1759_/B VGND VGND VPWR VPWR _2581_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1691_ _2391_/Q _2388_/Q VGND VGND VPWR VPWR _1693_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _2324_/A VGND VGND VPWR VPWR _2317_/A sky130_fd_sc_hd__buf_2
XFILLER_3_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2236_/Y _2240_/Y _2242_/X VGND VGND VPWR VPWR _2243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2174_ _2497_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2174_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2414__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1958_ _1962_/A VGND VGND VPWR VPWR _1958_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1889_ _1913_/A VGND VGND VPWR VPWR _1894_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2564__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1992__A _1993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2328__A _2329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2047__B _2451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2063__A _2247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1526__A0 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2238__A _2238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2587__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1812_ _2599_/Q _2596_/Q VGND VGND VPWR VPWR _1815_/D sky130_fd_sc_hd__and2_1
XFILLER_160_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1743_ _1702_/X _2408_/Q _1741_/X _1742_/Y VGND VGND VPWR VPWR _1745_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1674_ _1674_/A _1674_/B VGND VGND VPWR VPWR _2384_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1517__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2226_ _2220_/Y _2203_/X _2225_/Y VGND VGND VPWR VPWR _2536_/D sky130_fd_sc_hd__o21ai_1
XFILLER_41_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2157_ _2151_/Y _2154_/Y _2156_/X VGND VGND VPWR VPWR _2157_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ _2082_/Y _2071_/X _2087_/Y VGND VGND VPWR VPWR _2520_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__1987__A _1987_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1508__A0 _2450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1897__A _1900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1211__A2 _1191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1390_ _1390_/A VGND VGND VPWR VPWR _2504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1657__A1_N _1647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2011_ _2011_/A VGND VGND VPWR VPWR _2011_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1726_ _1722_/X _1727_/C _1727_/D _1727_/B VGND VGND VPWR VPWR _1728_/A sky130_fd_sc_hd__o22a_1
XFILLER_208_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1657_ _1647_/X _2420_/Q _1655_/X _1656_/Y VGND VGND VPWR VPWR _1660_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_208_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1588_ _1588_/A _2440_/Q _2443_/Q _2442_/Q VGND VGND VPWR VPWR _1588_/X sky130_fd_sc_hd__or4_1
XFILLER_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2053__C_N _2411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2209_ _2501_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2209_/X sky130_fd_sc_hd__o31a_1
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2028__D _2028_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2560_ _2560_/CLK _2560_/D _2317_/Y VGND VGND VPWR VPWR _2560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1196__A1 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1511_ _1511_/A VGND VGND VPWR VPWR _2449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2491_ _2560_/CLK _2491_/D _1986_/Y VGND VGND VPWR VPWR _2491_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1442_ _1486_/A VGND VGND VPWR VPWR _1451_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1373_ _1373_/A VGND VGND VPWR VPWR _2511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1671__A2 _1673_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1330__A _1374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1709_ _2397_/Q _2394_/Q VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__and2_1
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2071__A _2116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input67_A wbs_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2246__A _2246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1991_ _1993_/A VGND VGND VPWR VPWR _1991_/Y sky130_fd_sc_hd__inv_2
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _2569_/CLK _2543_/D VGND VGND VPWR VPWR _2543_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2474_ _2595_/CLK _2474_/D _1965_/Y VGND VGND VPWR VPWR _2474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1425_ _1425_/A VGND VGND VPWR VPWR _2488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1325__A _2170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1356_ input57/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1356_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ input41/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1995__A _1999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1235__A _2026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2066__A _2066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2470__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1210_ _1199_/Y _1207_/X _1209_/X _2577_/Q VGND VGND VPWR VPWR _2576_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2190_ _2499_/Q _2155_/X _2165_/X _2189_/X VGND VGND VPWR VPWR _2190_/X sky130_fd_sc_hd__o31a_1
XFILLER_211_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2264__C_N _2435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ _1974_/A VGND VGND VPWR VPWR _1974_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2051__A2 _2022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2526_ _2560_/CLK _2526_/D VGND VGND VPWR VPWR _2526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2457_ _2459_/CLK _2457_/D _1943_/Y VGND VGND VPWR VPWR _2457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1408_ _1430_/A VGND VGND VPWR VPWR _1417_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2388_ _2459_/CLK _2388_/D _1859_/Y VGND VGND VPWR VPWR _2388_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1339_ _1339_/A VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__buf_2
XFILLER_186_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2493__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2290__A2 _2116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2281__A2 _2066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2033__A2 _2074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ _2391_/Q _2388_/Q VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__and2_1
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1574__S _1578_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2311_/A VGND VGND VPWR VPWR _2311_/Y sky130_fd_sc_hd__inv_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2242_ _2505_/Q _2241_/X _2208_/X _2231_/X VGND VGND VPWR VPWR _2242_/X sky130_fd_sc_hd__o31a_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2173_ _1628_/C _2118_/X _2162_/X _2172_/Y VGND VGND VPWR VPWR _2173_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ _1975_/A VGND VGND VPWR VPWR _1962_/A sky130_fd_sc_hd__buf_2
XFILLER_198_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1888_ _2361_/A VGND VGND VPWR VPWR _1913_/A sky130_fd_sc_hd__buf_2
XFILLER_200_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2509_ _2512_/CLK _2509_/D _2008_/Y VGND VGND VPWR VPWR _2509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__A _2186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1732__A2_N _2409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1462__A0 _2471_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1811_ _2428_/Q VGND VGND VPWR VPWR _1815_/C sky130_fd_sc_hd__inv_2
XFILLER_19_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1742_ _2407_/Q _2402_/Q VGND VGND VPWR VPWR _1742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1673_ _1777_/A _1673_/B _1673_/C _1673_/D VGND VGND VPWR VPWR _1674_/B sky130_fd_sc_hd__nor4_1
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1517__A1 _2438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2221_/Y _2223_/Y _2224_/X VGND VGND VPWR VPWR _2225_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2156_ _2495_/Q _2155_/X _2122_/X _2146_/X VGND VGND VPWR VPWR _2156_/X sky130_fd_sc_hd__o31a_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2087_ _2083_/Y _2085_/Y _2086_/X VGND VGND VPWR VPWR _2087_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2531__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1508__A1 _2451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2074__A _2074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2404__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2249__A _2249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2010_ _2011_/A VGND VGND VPWR VPWR _2010_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2554__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1725_ _2401_/Q _2398_/Q VGND VGND VPWR VPWR _1727_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1656_ _2381_/Q _2378_/Q VGND VGND VPWR VPWR _1656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1587_ _2441_/Q VGND VGND VPWR VPWR _1588_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2208_ _2252_/A VGND VGND VPWR VPWR _2208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1998__A _1999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2139_ _2134_/Y _2137_/Y _2138_/X VGND VGND VPWR VPWR _2139_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2427__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A wbs_adr_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1196__A2 _1191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1510_ _2449_/Q _2450_/Q _1589_/A VGND VGND VPWR VPWR _1511_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2490_ _2512_/CLK _2490_/D _1985_/Y VGND VGND VPWR VPWR _2490_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1441_ _2448_/Q VGND VGND VPWR VPWR _1486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1372_ _2511_/Q _2512_/Q _1372_/S VGND VGND VPWR VPWR _1373_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2161__B _2161_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1708_ _2395_/Q _2392_/Q _1707_/B VGND VGND VPWR VPWR _2395_/D sky130_fd_sc_hd__a21o_1
XFILLER_69_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1639_ _2422_/Q VGND VGND VPWR VPWR _1643_/C sky130_fd_sc_hd__inv_2
XFILLER_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input4_A wbs_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ _1993_/A VGND VGND VPWR VPWR _1990_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ _2569_/CLK _2542_/D VGND VGND VPWR VPWR _2542_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2473_ _2595_/CLK _2473_/D _1964_/Y VGND VGND VPWR VPWR _2473_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1424_ _2488_/Q _2489_/Q _1428_/S VGND VGND VPWR VPWR _1425_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1355_ _1497_/A VGND VGND VPWR VPWR _1372_/S sky130_fd_sc_hd__buf_2
XFILLER_60_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1608_/B VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1341__A _2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1487__S _1495_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1251__A _1497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1323__A2 _1311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1973_ _1974_/A VGND VGND VPWR VPWR _1973_/Y sky130_fd_sc_hd__inv_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2525_ _2560_/CLK _2525_/D VGND VGND VPWR VPWR _2525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2456_ _2459_/CLK _2456_/D _1942_/Y VGND VGND VPWR VPWR _2456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1407_ _1407_/A VGND VGND VPWR VPWR _2496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2387_ _2459_/CLK _2387_/D _1856_/Y VGND VGND VPWR VPWR _2387_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1338_ _2553_/Q _1311_/X _1335_/X _1337_/Y VGND VGND VPWR VPWR _2552_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1269_ _2565_/Q VGND VGND VPWR VPWR _1269_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2042__A3 _2016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1246__A _1297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2077__A _2252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1241__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2311_/A VGND VGND VPWR VPWR _2310_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2241_/A VGND VGND VPWR VPWR _2241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2172_ _2187_/A _2465_/Q VGND VGND VPWR VPWR _2172_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1956_ _1956_/A VGND VGND VPWR VPWR _1956_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1887_ _1887_/A VGND VGND VPWR VPWR _1887_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2508_ _2512_/CLK _2508_/D _2007_/Y VGND VGND VPWR VPWR _2508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2460__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2439_ _2577_/CLK _2439_/D _1922_/Y VGND VGND VPWR VPWR _2439_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input42_A wbs_dat_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1810_ _2597_/Q _2594_/Q _1809_/B VGND VGND VPWR VPWR _2597_/D sky130_fd_sc_hd__a21o_1
XFILLER_73_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1741_ _2407_/Q _2402_/Q VGND VGND VPWR VPWR _1741_/X sky130_fd_sc_hd__and2_1
XFILLER_89_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2270__A _2542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1672_ _1672_/A VGND VGND VPWR VPWR _1777_/A sky130_fd_sc_hd__buf_2
XFILLER_201_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2483__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2503_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2224_/X sky130_fd_sc_hd__o31a_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2155_ _2241_/A VGND VGND VPWR VPWR _2155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2086_ _2487_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2086_/X sky130_fd_sc_hd__o31a_1
XFILLER_78_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1495__S _1495_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1939_ _1943_/A VGND VGND VPWR VPWR _1939_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2355__A _2355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2090__A _2170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2265__A _2272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1738__A2 _2439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1724_ _2401_/Q _2398_/Q VGND VGND VPWR VPWR _1727_/D sky130_fd_sc_hd__and2_1
XFILLER_69_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1655_ _2381_/Q _2378_/Q VGND VGND VPWR VPWR _1655_/X sky130_fd_sc_hd__and2_1
XFILLER_208_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1586_ _2445_/Q _1586_/B _2447_/Q _2446_/Q VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__or4b_1
XFILLER_99_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2207_ _1815_/C _2186_/X _2205_/X _2206_/Y VGND VGND VPWR VPWR _2207_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2379__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _2493_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2138_/X sky130_fd_sc_hd__o31a_1
XFILLER_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2069_ _2060_/Y _2022_/X _2068_/Y VGND VGND VPWR VPWR _2518_/D sky130_fd_sc_hd__o21ai_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2154__A2 _2118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1440_ _1440_/A VGND VGND VPWR VPWR _2481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2145__A2 _2135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1371_ _1371_/A VGND VGND VPWR VPWR _2512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2521__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1164__A _1200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1339__A _1339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1707_ _1707_/A _1707_/B VGND VGND VPWR VPWR _2394_/D sky130_fd_sc_hd__nor2_1
XFILLER_195_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1638_ _2375_/Q _2372_/Q _1637_/B VGND VGND VPWR VPWR _2375_/D sky130_fd_sc_hd__a21o_1
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1569_ _2186_/A VGND VGND VPWR VPWR _1578_/S sky130_fd_sc_hd__buf_2
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1583__A0 input35/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2544__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1712__A _1747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2541_ _2569_/CLK _2541_/D VGND VGND VPWR VPWR _2541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1574__A0 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2472_ _2595_/CLK _2472_/D _1962_/Y VGND VGND VPWR VPWR _2472_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1423_ _1423_/A VGND VGND VPWR VPWR _2489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1354_ _2550_/Q _1339_/X _1351_/X _1353_/Y VGND VGND VPWR VPWR _2549_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1285_ _2563_/Q _1261_/X _1282_/X _1284_/Y VGND VGND VPWR VPWR _2562_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2417__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2567__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1556__A0 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2257__B _2292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ _1974_/A VGND VGND VPWR VPWR _1972_/Y sky130_fd_sc_hd__inv_2
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2524_ _2560_/CLK _2524_/D VGND VGND VPWR VPWR _2524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2455_ _2459_/CLK _2455_/D _1941_/Y VGND VGND VPWR VPWR _2455_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1406_ _2496_/Q _2497_/Q _1406_/S VGND VGND VPWR VPWR _1407_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2386_ _2601_/CLK _2386_/D _1855_/Y VGND VGND VPWR VPWR _2386_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1337_ _1320_/X _1313_/X _1336_/Y VGND VGND VPWR VPWR _1337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1268_ _1293_/A VGND VGND VPWR VPWR _1268_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1199_ input58/X _1191_/X _1339_/A VGND VGND VPWR VPWR _1199_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_129_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1498__S _1506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2240_ _1243_/Y _2237_/X _2205_/X _2239_/Y VGND VGND VPWR VPWR _2240_/Y sky130_fd_sc_hd__o211ai_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2171_ _2171_/A _2228_/B VGND VGND VPWR VPWR _2171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1900__A _1900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1955_ _1956_/A VGND VGND VPWR VPWR _1955_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1886_ _1887_/A VGND VGND VPWR VPWR _1886_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2507_ _2576_/CLK _2507_/D _2005_/Y VGND VGND VPWR VPWR _2507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2438_ _2577_/CLK _2438_/D _1921_/Y VGND VGND VPWR VPWR _2438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2369_ _2599_/CLK _2369_/D _1835_/Y VGND VGND VPWR VPWR _2369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1220__B1_N _1339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input35_A wbs_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1740_ _1740_/A VGND VGND VPWR VPWR _2404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1671_ _1631_/X _1673_/C _1673_/D _1673_/B VGND VGND VPWR VPWR _1674_/A sky130_fd_sc_hd__o22a_1
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2223_ _1254_/Y _2135_/X _2205_/X _2222_/Y VGND VGND VPWR VPWR _2223_/Y sky130_fd_sc_hd__o211ai_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2154_ _1643_/C _2118_/X _2119_/X _2153_/Y VGND VGND VPWR VPWR _2154_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_187_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2085_ _1336_/Y _2062_/X _2074_/X _2084_/Y VGND VGND VPWR VPWR _2085_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1938_ _1944_/A VGND VGND VPWR VPWR _1943_/A sky130_fd_sc_hd__buf_2
XFILLER_33_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1869_ _1869_/A VGND VGND VPWR VPWR _1869_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2450__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1199__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1723_ _2410_/Q VGND VGND VPWR VPWR _1727_/C sky130_fd_sc_hd__clkinv_2
XFILLER_121_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1654_ _2379_/Q _2376_/Q _1653_/B VGND VGND VPWR VPWR _2379_/D sky130_fd_sc_hd__a21o_1
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1585_ _2444_/Q VGND VGND VPWR VPWR _1586_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2229_/A _2469_/Q VGND VGND VPWR VPWR _2206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2137_ _1304_/Y _2135_/X _2119_/X _2136_/Y VGND VGND VPWR VPWR _2137_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2068_ _2061_/Y _2065_/Y _2067_/X VGND VGND VPWR VPWR _2068_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_39_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2473__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1370_ _2512_/Q _2406_/Q _1372_/S VGND VGND VPWR VPWR _1371_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2081__A2 _2071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1706_ _1703_/X _1704_/Y _1706_/C _2413_/Q VGND VGND VPWR VPWR _1707_/B sky130_fd_sc_hd__and4bb_1
XFILLER_69_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1637_ _1637_/A _1637_/B VGND VGND VPWR VPWR _2374_/D sky130_fd_sc_hd__nor2_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1355__A _1497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1568_ _1568_/A VGND VGND VPWR VPWR _2415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1499_ _1499_/A VGND VGND VPWR VPWR _2455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2496__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2186__A _2186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1583__A1 _2408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1335__A1 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2369__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2540_ _2569_/CLK _2540_/D VGND VGND VPWR VPWR _2540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1169__B_N _2012_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2471_ _2595_/CLK _2471_/D _1961_/Y VGND VGND VPWR VPWR _2471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1422_ _2489_/Q _2490_/Q _1428_/S VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1353_ _1346_/X _1341_/X _1352_/Y VGND VGND VPWR VPWR _1353_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1284_ _1268_/X _1263_/X _2171_/A VGND VGND VPWR VPWR _1284_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2511__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input65_A wbs_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ _1974_/A VGND VGND VPWR VPWR _1971_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1795__A1 _1722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2523_ _2560_/CLK _2523_/D VGND VGND VPWR VPWR _2523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2454_ _2549_/CLK _2454_/D _1940_/Y VGND VGND VPWR VPWR _2454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1405_ _1405_/A VGND VGND VPWR VPWR _2497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2385_ _2601_/CLK _2385_/D _1854_/Y VGND VGND VPWR VPWR _2385_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1336_ _2552_/Q VGND VGND VPWR VPWR _1336_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 wb_rst_i VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
XFILLER_211_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1267_ input45/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1267_/X sky130_fd_sc_hd__o21ba_1
XFILLER_84_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1198_ _1497_/A VGND VGND VPWR VPWR _1339_/A sky130_fd_sc_hd__buf_2
XFILLER_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2534__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2170_ _2170_/A VGND VGND VPWR VPWR _2228_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2557__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1465__A0 _2470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2284__A _2544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1954_ _1956_/A VGND VGND VPWR VPWR _1954_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1885_ _1887_/A VGND VGND VPWR VPWR _1885_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1628__A _1643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2506_ _2576_/CLK _2506_/D _2004_/Y VGND VGND VPWR VPWR _2506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2437_ _2577_/CLK _2437_/D _1918_/Y VGND VGND VPWR VPWR _2437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2178__B _2228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2368_ _2599_/CLK _2368_/D _1834_/Y VGND VGND VPWR VPWR _2368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ _2066_/A VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2299_ input1/X VGND VGND VPWR VPWR _2324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2194__A _2194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input28_A wbs_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1447__A0 _2478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1670_ _2385_/Q _2382_/Q VGND VGND VPWR VPWR _1673_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__A _2294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1183__A _1183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2222_ _2229_/A _2471_/Q VGND VGND VPWR VPWR _2222_/Y sky130_fd_sc_hd__nand2_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2153_ _2187_/A _2463_/Q VGND VGND VPWR VPWR _2153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1911__A _1912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2084_ _2099_/A _2455_/Q VGND VGND VPWR VPWR _2084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1937_ _1937_/A VGND VGND VPWR VPWR _1937_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1868_ _1869_/A VGND VGND VPWR VPWR _1868_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1799_ _2595_/Q _2592_/Q VGND VGND VPWR VPWR _1799_/X sky130_fd_sc_hd__and2_1
XFILLER_176_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2189__A _2231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2560_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2099__A _2099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2093__B1 _2074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1199__A2 _1191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1178__A _1178_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1722_ _1722_/A VGND VGND VPWR VPWR _1722_/X sky130_fd_sc_hd__buf_2
XFILLER_34_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1653_ _1653_/A _1653_/B VGND VGND VPWR VPWR _2378_/D sky130_fd_sc_hd__nor2_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1584_ _1584_/A VGND VGND VPWR VPWR _2408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2249_/A VGND VGND VPWR VPWR _2205_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2136_ _2144_/A _2461_/Q VGND VGND VPWR VPWR _2136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1234__B1_N _1224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2067_ _2485_/Q _2066_/X _2016_/X _2056_/X VGND VGND VPWR VPWR _2067_/X sky130_fd_sc_hd__o31a_1
XFILLER_54_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1705_ _1702_/X _2413_/Q _1703_/X _1704_/Y VGND VGND VPWR VPWR _1707_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1636__A _1643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1636_ _1643_/A _1636_/B _1636_/C _1636_/D VGND VGND VPWR VPWR _1637_/B sky130_fd_sc_hd__nor4_1
XFILLER_86_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1567_ input64/X _2415_/Q _1567_/S VGND VGND VPWR VPWR _1568_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1344__A2 _1339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1498_ _2455_/Q _2456_/Q _1506_/S VGND VGND VPWR VPWR _1499_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2119_ _2249_/A VGND VGND VPWR VPWR _2119_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2440__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2296__B1 _2032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input10_A wbs_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2590__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _2595_/CLK _2470_/D _1960_/Y VGND VGND VPWR VPWR _2470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1421_ _1421_/A VGND VGND VPWR VPWR _2490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1352_ _2549_/Q VGND VGND VPWR VPWR _1352_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1283_ _2562_/Q VGND VGND VPWR VPWR _2171_/A sky130_fd_sc_hd__inv_2
XFILLER_81_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1191__A _2237_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2287__B1 _2074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2463__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1619_ _2371_/Q _2368_/Q VGND VGND VPWR VPWR _1621_/B sky130_fd_sc_hd__nor2_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2599_ _2599_/CLK _2599_/D _2365_/Y VGND VGND VPWR VPWR _2599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A wbs_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1253__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input58_A wbs_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ _1974_/A VGND VGND VPWR VPWR _1970_/Y sky130_fd_sc_hd__inv_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2486__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1186__A input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2522_ _2553_/CLK _2522_/D VGND VGND VPWR VPWR _2522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2453_ _2459_/CLK _2453_/D _1939_/Y VGND VGND VPWR VPWR _2453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1404_ _2497_/Q _2498_/Q _1406_/S VGND VGND VPWR VPWR _1405_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2384_ _2601_/CLK _2384_/D _1853_/Y VGND VGND VPWR VPWR _2384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1335_ input63/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1335_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 wbs_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
X_1266_ _2567_/Q _1261_/X _1262_/X _1265_/Y VGND VGND VPWR VPWR _2566_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1197_ _2448_/Q VGND VGND VPWR VPWR _1497_/A sky130_fd_sc_hd__buf_2
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2561__RESET_B _2319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1465__A1 _2471_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1953_ _1956_/A VGND VGND VPWR VPWR _1953_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1909__A _1912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1884_ _1887_/A VGND VGND VPWR VPWR _1884_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2505_ _2512_/CLK _2505_/D _2003_/Y VGND VGND VPWR VPWR _2505_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2436_ _2577_/CLK _2436_/D _1917_/Y VGND VGND VPWR VPWR _2436_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2367_ _2367_/A VGND VGND VPWR VPWR _2367_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2501__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1318_ _1512_/D VGND VGND VPWR VPWR _2066_/A sky130_fd_sc_hd__buf_2
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2298_ _2291_/Y _2116_/A _2297_/Y VGND VGND VPWR VPWR _2545_/D sky130_fd_sc_hd__o21ai_2
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1249_ _1242_/X _1237_/X _2228_/A VGND VGND VPWR VPWR _1249_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2194__B _2236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output89_A _2541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2524__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__B _2478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1183__B input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2221_ _2264_/A _2236_/B _2430_/Q VGND VGND VPWR VPWR _2221_/Y sky130_fd_sc_hd__nor3b_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2152_ _2238_/A VGND VGND VPWR VPWR _2187_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2083_ _2083_/A _2134_/B _2414_/Q VGND VGND VPWR VPWR _2083_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1936_ _1937_/A VGND VGND VPWR VPWR _1936_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1867_ _1869_/A VGND VGND VPWR VPWR _1867_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput60 wbs_dat_i[3] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_2
XFILLER_50_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1798_ _2593_/Q _2590_/Q _1797_/B VGND VGND VPWR VPWR _2593_/D sky130_fd_sc_hd__a21o_1
XFILLER_85_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1374__A _1374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2419_ _2560_/CLK _2419_/D _1897_/Y VGND VGND VPWR VPWR _2419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2547__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input40_A wbs_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1721_ _2399_/Q _2396_/Q _1720_/B VGND VGND VPWR VPWR _2399_/D sky130_fd_sc_hd__a21o_1
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1652_ _1648_/X _1649_/Y _1652_/C _2421_/Q VGND VGND VPWR VPWR _1653_/B sky130_fd_sc_hd__and4bb_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1583_ input35/X _2408_/Q _1583_/S VGND VGND VPWR VPWR _1584_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1194__A _1589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2204_ _2204_/A _2228_/B VGND VGND VPWR VPWR _2204_/Y sky130_fd_sc_hd__nor2_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2135_ _2237_/A VGND VGND VPWR VPWR _2135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2066_ _2066_/A VGND VGND VPWR VPWR _2066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1919_ _2361_/A VGND VGND VPWR VPWR _1944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1832__A _2361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1356__B1_N _1372_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2292__B _2292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1189__A _2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1704_ _2395_/Q _2392_/Q VGND VGND VPWR VPWR _1704_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ _1631_/X _1636_/C _1636_/D _1636_/B VGND VGND VPWR VPWR _1637_/A sky130_fd_sc_hd__o22a_1
XFILLER_144_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1566_ _1566_/A VGND VGND VPWR VPWR _2416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1497_ _1497_/A VGND VGND VPWR VPWR _1506_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_113_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ _2186_/A VGND VGND VPWR VPWR _2118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2049_ _2483_/Q _1346_/A _2016_/X _2246_/A VGND VGND VPWR VPWR _2049_/X sky130_fd_sc_hd__o31a_1
XFILLER_93_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2048__A1 _1727_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1420_ _2490_/Q _2491_/Q _1428_/S VGND VGND VPWR VPWR _1421_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1351_ input60/X _2046_/B _1330_/X VGND VGND VPWR VPWR _1351_/X sky130_fd_sc_hd__o21ba_1
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1282_ input42/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__o21ba_1
XFILLER_205_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1647__A _1747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1618_ _2371_/Q _2368_/Q VGND VGND VPWR VPWR _1621_/D sky130_fd_sc_hd__and2_1
XFILLER_138_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2598_ _2599_/CLK _2598_/D _2364_/Y VGND VGND VPWR VPWR _2598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1549_ _1549_/A VGND VGND VPWR VPWR _2424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2521_ _2553_/CLK _2521_/D VGND VGND VPWR VPWR _2521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2452_ _2549_/CLK _2452_/D _1937_/Y VGND VGND VPWR VPWR _2452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1403_ _1403_/A VGND VGND VPWR VPWR _2498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2383_ _2601_/CLK _2383_/D _1852_/Y VGND VGND VPWR VPWR _2383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1334_ _2554_/Q _1311_/X _1331_/X _1333_/Y VGND VGND VPWR VPWR _2553_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1265_ _1242_/X _1263_/X _2204_/A VGND VGND VPWR VPWR _1265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput3 wbs_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1196_ input59/X _1191_/X _1195_/Y VGND VGND VPWR VPWR _2577_/D sky130_fd_sc_hd__o21a_1
XFILLER_149_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2580__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2001__A _2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _1956_/A VGND VGND VPWR VPWR _1952_/Y sky130_fd_sc_hd__inv_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1883_ _1887_/A VGND VGND VPWR VPWR _1883_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1197__A _2448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2504_ _2576_/CLK _2504_/D _2002_/Y VGND VGND VPWR VPWR _2504_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2435_ _2577_/CLK _2435_/D _1916_/Y VGND VGND VPWR VPWR _2435_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2366_ _2366_/A VGND VGND VPWR VPWR _2366_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1317_ input66/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1317_/X sky130_fd_sc_hd__o21ba_1
XFILLER_22_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2297_ _2292_/Y _2295_/Y _2296_/X VGND VGND VPWR VPWR _2297_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1248_ _2569_/Q VGND VGND VPWR VPWR _2228_/A sky130_fd_sc_hd__inv_2
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1179_ _1179_/A input2/X VGND VGND VPWR VPWR _1182_/A sky130_fd_sc_hd__nor2_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2476__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2536_/Q VGND VGND VPWR VPWR _2220_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2151_ _2151_/A _2161_/B VGND VGND VPWR VPWR _2151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2082_ _2520_/Q VGND VGND VPWR VPWR _2082_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1935_ _1937_/A VGND VGND VPWR VPWR _1935_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1866_ _1869_/A VGND VGND VPWR VPWR _1866_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1743__A2_N _2408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput50 wbs_dat_i[23] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput61 wbs_dat_i[4] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1797_ _1797_/A _1797_/B VGND VGND VPWR VPWR _2592_/D sky130_fd_sc_hd__nor2_1
XFILLER_190_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2418_ _2560_/CLK _2418_/D _1896_/Y VGND VGND VPWR VPWR _2418_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2499__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2349_ _2355_/A VGND VGND VPWR VPWR _2354_/A sky130_fd_sc_hd__buf_2
XFILLER_131_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input33_A wbs_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1504__S _1506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2093__A2 _1583_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1720_ _1720_/A _1720_/B VGND VGND VPWR VPWR _2398_/D sky130_fd_sc_hd__nor2_1
XFILLER_160_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1651_ _2546_/Q VGND VGND VPWR VPWR _1652_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_176_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1582_ _1582_/A VGND VGND VPWR VPWR _2409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1356__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2203_ _2246_/A VGND VGND VPWR VPWR _2203_/X sky130_fd_sc_hd__clkbuf_2
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2134_ _2194_/A _2134_/B _2420_/Q VGND VGND VPWR VPWR _2134_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_67_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2065_ _1347_/Y _2062_/X _2030_/X _2064_/Y VGND VGND VPWR VPWR _2065_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_78_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1918_ _1918_/A VGND VGND VPWR VPWR _1918_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1849_ _1850_/A VGND VGND VPWR VPWR _1849_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1385__A _2448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2514__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1510__A1 _2450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1189__B _1512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1703_ _2395_/Q _2392_/Q VGND VGND VPWR VPWR _1703_/X sky130_fd_sc_hd__and2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1634_ _2375_/Q _2372_/Q VGND VGND VPWR VPWR _1636_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1565_ input65/X _2416_/Q _1567_/S VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1496_ _1496_/A VGND VGND VPWR VPWR _2456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2537__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2117_ _2117_/A _2161_/B VGND VGND VPWR VPWR _2117_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2048_ _1727_/C _1583_/S _2030_/X _2047_/Y VGND VGND VPWR VPWR _2048_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_58_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2004__A _2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2296__A2 _2066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2048__A2 _1583_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1737__B _2439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1350_ _2170_/A VGND VGND VPWR VPWR _2046_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1281_ _2564_/Q _1261_/X _1278_/X _1280_/Y VGND VGND VPWR VPWR _2563_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2287__A2 _1297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1617_ _2425_/Q VGND VGND VPWR VPWR _1621_/C sky130_fd_sc_hd__inv_2
XFILLER_47_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2597_ _2599_/CLK _2597_/D _2363_/Y VGND VGND VPWR VPWR _2597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1548_ input42/X _2424_/Q _1556_/S VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1479_ _1479_/A VGND VGND VPWR VPWR _2464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2269__A2 _2246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2520_ _2553_/CLK _2520_/D VGND VGND VPWR VPWR _2520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2451_ _2549_/CLK _2451_/D _1936_/Y VGND VGND VPWR VPWR _2451_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ _2498_/Q _2499_/Q _1406_/S VGND VGND VPWR VPWR _1403_/A sky130_fd_sc_hd__mux2_1
X_2382_ _2459_/CLK _2382_/D _1850_/Y VGND VGND VPWR VPWR _2382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1333_ _1320_/X _1313_/X _2091_/A VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1264_ _2566_/Q VGND VGND VPWR VPWR _2204_/A sky130_fd_sc_hd__inv_2
XFILLER_83_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 wbs_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1195_ _2292_/A _1191_/X _1194_/X VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_168_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1658__A _1747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1247__B1_N _1224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input63_A wbs_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1951_ _1975_/A VGND VGND VPWR VPWR _1956_/A sky130_fd_sc_hd__buf_2
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1882_ _1882_/A VGND VGND VPWR VPWR _1887_/A sky130_fd_sc_hd__buf_2
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2503_ _2576_/CLK _2503_/D _2001_/Y VGND VGND VPWR VPWR _2503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2434_ _2577_/CLK _2434_/D _1915_/Y VGND VGND VPWR VPWR _2434_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2365_ _2366_/A VGND VGND VPWR VPWR _2365_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1316_ _2557_/Q _1311_/X _1312_/X _1315_/Y VGND VGND VPWR VPWR _2556_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2296_ _2512_/Q _2066_/A _2165_/A _2032_/X VGND VGND VPWR VPWR _2296_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1247_ input50/X _1246_/X _1224_/X VGND VGND VPWR VPWR _1247_/X sky130_fd_sc_hd__o21ba_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1178_ _1178_/A _1178_/B VGND VGND VPWR VPWR _2028_/B sky130_fd_sc_hd__nor2_8
XFILLER_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2012__A _2448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1604__B1 _1194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ _2528_/Q VGND VGND VPWR VPWR _2150_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2420__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2081_ _2070_/Y _2071_/X _2080_/Y VGND VGND VPWR VPWR _2519_/D sky130_fd_sc_hd__o21ai_1
XFILLER_4_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2570__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1934_ _1937_/A VGND VGND VPWR VPWR _1934_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1865_ _1869_/A VGND VGND VPWR VPWR _1865_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput40 wbs_dat_i[14] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput51 wbs_dat_i[24] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
Xinput62 wbs_dat_i[5] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_2
X_1796_ _1828_/A _1796_/B _1796_/C _1796_/D VGND VGND VPWR VPWR _1797_/B sky130_fd_sc_hd__nor4_1
XFILLER_122_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2417_ _2549_/CLK _2417_/D _1894_/Y VGND VGND VPWR VPWR _2417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2348_ _2348_/A VGND VGND VPWR VPWR _2348_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2279_ _2294_/A _2478_/Q VGND VGND VPWR VPWR _2279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2007__A _2011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2443__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input26_A wbs_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2593__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _1647_/X _2421_/Q _1648_/X _1649_/Y VGND VGND VPWR VPWR _1653_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output94_A _2545_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1581_ input46/X _2409_/Q _1583_/S VGND VGND VPWR VPWR _1582_/A sky130_fd_sc_hd__mux2_1
XFILLER_193_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2534_/Q VGND VGND VPWR VPWR _2202_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2133_ _2526_/Q VGND VGND VPWR VPWR _2133_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2064_ _2099_/A _2453_/Q VGND VGND VPWR VPWR _2064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1292__A1 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1917_ _1918_/A VGND VGND VPWR VPWR _1917_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1848_ _1850_/A VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2466__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1779_ _2587_/Q _2584_/Q _1778_/B VGND VGND VPWR VPWR _2587_/D sky130_fd_sc_hd__a21o_1
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1338__A2 _1311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1189__C _2028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2489__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2223__B1 _2205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1702_ _1747_/A VGND VGND VPWR VPWR _1702_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1633_ _2375_/Q _2372_/Q VGND VGND VPWR VPWR _1636_/D sky130_fd_sc_hd__and2_1
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1329__A2 _1311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1564_ _1564_/A VGND VGND VPWR VPWR _2417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1495_ _2456_/Q _2457_/Q _1495_/S VGND VGND VPWR VPWR _1496_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1652__C _1652_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2116_ _2116_/A VGND VGND VPWR VPWR _2116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2047_ _2054_/A _2451_/Q VGND VGND VPWR VPWR _2047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2057__A3 _2016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1820__A1_N _1652_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2020__A _2231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2601_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1280_ _1268_/X _1263_/X _2178_/A VGND VGND VPWR VPWR _1280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1247__A1 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1616_ _1672_/A VGND VGND VPWR VPWR _1828_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2596_ _2601_/CLK _2596_/D _2362_/Y VGND VGND VPWR VPWR _2596_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2504__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1547_ _1558_/A VGND VGND VPWR VPWR _1556_/S sky130_fd_sc_hd__buf_2
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1478_ _2464_/Q _2465_/Q _1484_/S VGND VGND VPWR VPWR _1479_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2015__A _2028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1229__A1 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2527__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2450_ _2549_/CLK _2450_/D _1935_/Y VGND VGND VPWR VPWR _2450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1401_ _1401_/A VGND VGND VPWR VPWR _2499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2381_ _2601_/CLK _2381_/D _1849_/Y VGND VGND VPWR VPWR _2381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1332_ _2553_/Q VGND VGND VPWR VPWR _2091_/A sky130_fd_sc_hd__inv_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1263_ _2024_/B VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 wbs_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1194_ _1589_/A VGND VGND VPWR VPWR _1194_/X sky130_fd_sc_hd__buf_4
XFILLER_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2579_ _2595_/CLK _2579_/D _2341_/Y VGND VGND VPWR VPWR _2579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input56_A wbs_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1950_ input1/X VGND VGND VPWR VPWR _1975_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1881_ _1881_/A VGND VGND VPWR VPWR _1881_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2502_ _2512_/CLK _2502_/D _1999_/Y VGND VGND VPWR VPWR _2502_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2433_ _2577_/CLK _2433_/D _1914_/Y VGND VGND VPWR VPWR _2433_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2364_ _2366_/A VGND VGND VPWR VPWR _2364_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1315_ _1293_/X _1313_/X _2117_/A VGND VGND VPWR VPWR _1315_/Y sky130_fd_sc_hd__o21ai_1
X_2295_ _2293_/Y _2186_/X _2074_/A _2294_/Y VGND VGND VPWR VPWR _2295_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1433__S _1439_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1246_ _1297_/A VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2102__A2 _2066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1177_ _1177_/A _1177_/B _1177_/C _1177_/D VGND VGND VPWR VPWR _1178_/B sky130_fd_sc_hd__nand4_4
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2012__B _2012_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2372__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__B1 _1643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2203__A _2246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2080_ _2073_/Y _2076_/Y _2079_/X VGND VGND VPWR VPWR _2080_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1933_ _1937_/A VGND VGND VPWR VPWR _1933_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1864_ _1882_/A VGND VGND VPWR VPWR _1869_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 wbs_adr_i[6] VGND VGND VPWR VPWR _1166_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput41 wbs_dat_i[15] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput52 wbs_dat_i[25] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput63 wbs_dat_i[6] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_2
X_1795_ _1722_/X _1796_/C _1796_/D _1796_/B VGND VGND VPWR VPWR _1797_/A sky130_fd_sc_hd__o22a_1
XFILLER_190_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2416_ _2560_/CLK _2416_/D _1893_/Y VGND VGND VPWR VPWR _2416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2347_ _2348_/A VGND VGND VPWR VPWR _2347_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2278_ _2285_/A _2285_/B _2437_/Q VGND VGND VPWR VPWR _2278_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_6_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1229_ input53/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1229_/X sky130_fd_sc_hd__o21ba_1
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2023__A _2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input19_A wbs_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1580_ _2186_/A VGND VGND VPWR VPWR _1583_/S sky130_fd_sc_hd__buf_2
XFILLER_67_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2193_/Y _2160_/X _2200_/Y VGND VGND VPWR VPWR _2533_/D sky130_fd_sc_hd__o21ai_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2132_ _2126_/Y _2116_/X _2131_/Y VGND VGND VPWR VPWR _2525_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2063_ _2247_/A VGND VGND VPWR VPWR _2099_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2108__A _2247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1916_ _1918_/A VGND VGND VPWR VPWR _1916_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1847_ _1850_/A VGND VGND VPWR VPWR _1847_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1778_ _1778_/A _1778_/B VGND VGND VPWR VPWR _2586_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1504__A0 _2452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2018__A _2514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1857__A _2361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2410__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2560__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1701_ _2393_/Q _2390_/Q _1700_/B VGND VGND VPWR VPWR _2393_/D sky130_fd_sc_hd__a21o_1
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1632_ _2423_/Q VGND VGND VPWR VPWR _1636_/C sky130_fd_sc_hd__inv_2
XFILLER_12_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1563_ input66/X _2417_/Q _1567_/S VGND VGND VPWR VPWR _1564_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1494_ _1494_/A VGND VGND VPWR VPWR _2457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2115_ _2524_/Q VGND VGND VPWR VPWR _2115_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2046_ _2046_/A _2046_/B VGND VGND VPWR VPWR _2046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_208_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2583__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2301__A _2305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1497__A _1497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1615_ _1615_/A VGND VGND VPWR VPWR _2447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2595_ _2595_/CLK _2595_/D _2360_/Y VGND VGND VPWR VPWR _2595_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1546_ _1546_/A VGND VGND VPWR VPWR _2425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1477_ _1477_/A VGND VGND VPWR VPWR _2465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _2249_/A VGND VGND VPWR VPWR _2074_/A sky130_fd_sc_hd__buf_2
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1200__A _1200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1756__A2_N _2437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2479__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2206__A _2229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1400_ _2499_/Q _2500_/Q _1406_/S VGND VGND VPWR VPWR _1401_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2380_ _2601_/CLK _2380_/D _1848_/Y VGND VGND VPWR VPWR _2380_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1331_ input64/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__o21ba_1
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1262_ input47/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__o21ba_1
XFILLER_211_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 wbs_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1193_ _2448_/Q VGND VGND VPWR VPWR _1589_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2116__A _2116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2578_ _2595_/CLK _2578_/D _2340_/Y VGND VGND VPWR VPWR _2578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1529_ _1529_/A VGND VGND VPWR VPWR _2433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2026__A _2026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input49_A wbs_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1880_ _1881_/A VGND VGND VPWR VPWR _1880_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2501_ _2576_/CLK _2501_/D _1998_/Y VGND VGND VPWR VPWR _2501_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2432_ _2577_/CLK _2432_/D _1912_/Y VGND VGND VPWR VPWR _2432_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2363_ _2366_/A VGND VGND VPWR VPWR _2363_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1314_ _2556_/Q VGND VGND VPWR VPWR _2117_/A sky130_fd_sc_hd__inv_2
XFILLER_135_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2294_ _2294_/A _2480_/Q VGND VGND VPWR VPWR _2294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1245_ _2571_/Q _1233_/X _1241_/X _1244_/Y VGND VGND VPWR VPWR _2570_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2102__A3 _2078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1176_ _1176_/A _1176_/B VGND VGND VPWR VPWR _1177_/D sky130_fd_sc_hd__nor2_2
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1788__A1_N _1652_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2517__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2096__A2 _2071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ _1944_/A VGND VGND VPWR VPWR _1937_/A sky130_fd_sc_hd__buf_2
XFILLER_128_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1863_ _1863_/A VGND VGND VPWR VPWR _1863_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput20 wbs_adr_i[26] VGND VGND VPWR VPWR _1176_/B sky130_fd_sc_hd__clkbuf_1
Xinput31 wbs_adr_i[7] VGND VGND VPWR VPWR _1166_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 wbs_dat_i[16] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
X_1794_ _2593_/Q _2590_/Q VGND VGND VPWR VPWR _1796_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput53 wbs_dat_i[26] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_2
Xinput64 wbs_dat_i[7] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2415_ _2560_/CLK _2415_/D _1892_/Y VGND VGND VPWR VPWR _2415_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2346_ _2348_/A VGND VGND VPWR VPWR _2346_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2277_ _2543_/Q VGND VGND VPWR VPWR _2277_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1228_ _2574_/Q _1209_/X _1225_/X _1227_/Y VGND VGND VPWR VPWR _2573_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2304__A _2305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1650__A1_N _1647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2214__A _2264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2200_ _2194_/Y _2197_/Y _2199_/X VGND VGND VPWR VPWR _2200_/Y sky130_fd_sc_hd__o21ai_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _2127_/Y _2129_/Y _2130_/X VGND VGND VPWR VPWR _2131_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2062_ _2170_/A VGND VGND VPWR VPWR _2062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2069__A2 _2022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ _1918_/A VGND VGND VPWR VPWR _1915_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1439__S _1439_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1846_ _1850_/A VGND VGND VPWR VPWR _1846_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1777_ _1777_/A _1777_/B _1777_/C _1777_/D VGND VGND VPWR VPWR _1778_/B sky130_fd_sc_hd__nor4_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1963__A _1975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2329_/A VGND VGND VPWR VPWR _2329_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1203__A _1512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input31_A wbs_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2223__A2 _2135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ _1700_/A _1700_/B VGND VGND VPWR VPWR _2392_/D sky130_fd_sc_hd__nor2_1
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1631_ _1672_/A VGND VGND VPWR VPWR _1631_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2385__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1562_ _1562_/A VGND VGND VPWR VPWR _2418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1493_ _2457_/Q _2458_/Q _1495_/S VGND VGND VPWR VPWR _1494_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2114_ _2105_/Y _2071_/X _2113_/Y VGND VGND VPWR VPWR _2523_/D sky130_fd_sc_hd__o21ai_1
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2045_ _2516_/Q VGND VGND VPWR VPWR _2045_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2119__A _2249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1829_ _1829_/A _1829_/B VGND VGND VPWR VPWR _2368_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1693__A _1777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2029__A _2249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1614_ _1614_/A _1614_/B _1614_/C VGND VGND VPWR VPWR _1615_/A sky130_fd_sc_hd__and3_1
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1199__B1_N _1339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2594_ _2599_/CLK _2594_/D _2359_/Y VGND VGND VPWR VPWR _2594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1545_ input43/X _2425_/Q _1545_/S VGND VGND VPWR VPWR _1546_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1476_ _2465_/Q _2466_/Q _1484_/S VGND VGND VPWR VPWR _1477_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2028_ _2213_/A _2028_/B _2028_/C _2028_/D VGND VGND VPWR VPWR _2249_/A sky130_fd_sc_hd__nand4_4
XFILLER_93_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2550__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2015__C _2028_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2312__A _2324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2222__A _2229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1330_ _1374_/A VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2423__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1261_ _1608_/B VGND VGND VPWR VPWR _1261_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1192_ _2577_/Q VGND VGND VPWR VPWR _2292_/A sky130_fd_sc_hd__inv_2
Xinput7 wbs_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2573__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2577_ _2577_/CLK _2577_/D _2339_/Y VGND VGND VPWR VPWR _2577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1528_ input52/X _2433_/Q _1534_/S VGND VGND VPWR VPWR _1529_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1459_ _1459_/A VGND VGND VPWR VPWR _2473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2446__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1881__A _1881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2596__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2500_ _2512_/CLK _2500_/D _1997_/Y VGND VGND VPWR VPWR _2500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2431_ _2569_/CLK _2431_/D _1911_/Y VGND VGND VPWR VPWR _2431_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2362_ _2366_/A VGND VGND VPWR VPWR _2362_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1313_ _2024_/B VGND VGND VPWR VPWR _1313_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2293_ _2439_/Q VGND VGND VPWR VPWR _2293_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1244_ _1242_/X _1237_/X _1243_/Y VGND VGND VPWR VPWR _1244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1175_ _1175_/A _1175_/B VGND VGND VPWR VPWR _1177_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2127__A _2194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2469__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2037__A _2285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2262__B1 _2261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__A2 _2061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input61_A wbs_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ _1931_/A VGND VGND VPWR VPWR _1931_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1862_ _1863_/A VGND VGND VPWR VPWR _1862_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput10 wbs_adr_i[17] VGND VGND VPWR VPWR _1183_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput21 wbs_adr_i[27] VGND VGND VPWR VPWR _1176_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput32 wbs_adr_i[8] VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__clkbuf_1
X_1793_ _2593_/Q _2590_/Q VGND VGND VPWR VPWR _1796_/D sky130_fd_sc_hd__and2_1
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput43 wbs_dat_i[17] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__A2 _1339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput54 wbs_dat_i[27] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_2
XFILLER_50_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput65 wbs_dat_i[8] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2414_ _2549_/CLK _2414_/D _1891_/Y VGND VGND VPWR VPWR _2414_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2345_ _2348_/A VGND VGND VPWR VPWR _2345_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2276_ _2270_/Y _2246_/X _2275_/Y VGND VGND VPWR VPWR _2542_/D sky130_fd_sc_hd__o21ai_1
XFILLER_42_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1227_ _1212_/X _1214_/X _1226_/Y VGND VGND VPWR VPWR _1227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2320__A _2323_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1370__S _1372_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2214__B _2236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2558__RESET_B _2315_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ _2492_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2130_/X sky130_fd_sc_hd__o31a_1
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2061_ _2083_/A _2061_/B _2412_/Q VGND VGND VPWR VPWR _2061_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_43_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1914_ _1918_/A VGND VGND VPWR VPWR _1914_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1845_ _2367_/A VGND VGND VPWR VPWR _1850_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1776_ _1722_/X _1777_/C _1777_/D _1777_/B VGND VGND VPWR VPWR _1778_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2507__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2329_/A VGND VGND VPWR VPWR _2328_/Y sky130_fd_sc_hd__inv_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2259_ _1777_/C _2186_/X _2249_/X _2258_/Y VGND VGND VPWR VPWR _2259_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_211_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1203__B _2028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2315__A _2317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A wbs_adr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1630_ _2373_/Q _2370_/Q _1629_/B VGND VGND VPWR VPWR _2373_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output92_A _2516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1561_ input36/X _2418_/Q _1567_/S VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1195__B1 _1194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1492_ _1492_/A VGND VGND VPWR VPWR _2458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2113_ _2107_/Y _2110_/Y _2112_/X VGND VGND VPWR VPWR _2113_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2044_ _2036_/Y _2022_/X _2043_/Y VGND VGND VPWR VPWR _2515_/D sky130_fd_sc_hd__o21ai_1
XFILLER_110_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2135__A _2237_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1664__A1_N _1647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1828_ _1828_/A _1828_/B _1828_/C _1828_/D VGND VGND VPWR VPWR _1829_/B sky130_fd_sc_hd__nor4_1
XFILLER_30_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1759_ _1759_/A _1759_/B VGND VGND VPWR VPWR _2580_/D sky130_fd_sc_hd__nor2_1
XFILLER_190_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1214__A _2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2045__A _2516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1613_ _2445_/Q _1586_/B _2446_/Q _1606_/C _2447_/Q VGND VGND VPWR VPWR _1614_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_103_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2593_ _2599_/CLK _2593_/D _2358_/Y VGND VGND VPWR VPWR _2593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1544_ _1544_/A VGND VGND VPWR VPWR _2426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1475_ _1486_/A VGND VGND VPWR VPWR _1484_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_141_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1969__A _1975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2027_ _2294_/A _2449_/Q VGND VGND VPWR VPWR _2027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1209__A _1608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1879__A _1881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2375__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1764__D _2436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2222__B _2471_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1570__A0 input63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1260_ _2568_/Q _1233_/X _1257_/X _1259_/Y VGND VGND VPWR VPWR _2567_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2114__A2 _2071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1191_ _2237_/A VGND VGND VPWR VPWR _1191_/X sky130_fd_sc_hd__clkbuf_4
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 wbs_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2576_ _2576_/CLK _2576_/D _2338_/Y VGND VGND VPWR VPWR _2576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1527_ _1527_/A VGND VGND VPWR VPWR _2434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1458_ _2473_/Q _2474_/Q _1462_/S VGND VGND VPWR VPWR _1459_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1389_ _2504_/Q _2505_/Q _1395_/S VGND VGND VPWR VPWR _1390_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2323__A _2323_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1552__A0 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2430_ _2577_/CLK _2430_/D _1910_/Y VGND VGND VPWR VPWR _2430_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2361_ _2361_/A VGND VGND VPWR VPWR _2366_/A sky130_fd_sc_hd__buf_2
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2540__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1312_ input36/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1312_/X sky130_fd_sc_hd__o21ba_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2292_ _2292_/A _2292_/B VGND VGND VPWR VPWR _2292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1243_ _2570_/Q VGND VGND VPWR VPWR _1243_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1174_ _1174_/A _1174_/B VGND VGND VPWR VPWR _1177_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2127__B _2134_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2143__A _2194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1982__A _2006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2559_ _2560_/CLK _2559_/D _2316_/Y VGND VGND VPWR VPWR _2559_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1534__A0 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2318__A _2324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2413__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2053__A _2083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1892__A _1894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2563__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_A wbs_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1931_/A VGND VGND VPWR VPWR _1930_/Y sky130_fd_sc_hd__inv_2
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1861_ _1863_/A VGND VGND VPWR VPWR _1861_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 wbs_adr_i[18] VGND VGND VPWR VPWR _1184_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 wbs_adr_i[28] VGND VGND VPWR VPWR _1172_/B sky130_fd_sc_hd__clkbuf_1
X_1792_ _2431_/Q VGND VGND VPWR VPWR _1796_/C sky130_fd_sc_hd__inv_2
Xinput33 wbs_adr_i[9] VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput44 wbs_dat_i[18] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput55 wbs_dat_i[28] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput66 wbs_dat_i[9] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2413_ _2549_/CLK _2413_/D _1890_/Y VGND VGND VPWR VPWR _2413_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2344_ _2348_/A VGND VGND VPWR VPWR _2344_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2275_ _2271_/Y _2273_/Y _2274_/X VGND VGND VPWR VPWR _2275_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_6_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1226_ _2573_/Q VGND VGND VPWR VPWR _1226_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1977__A _1980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2586__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1561__S _1567_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2060_ _2518_/Q VGND VGND VPWR VPWR _2060_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1769__A2_N _2435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A VGND VGND VPWR VPWR _1918_/A sky130_fd_sc_hd__buf_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1844_ _1844_/A VGND VGND VPWR VPWR _1844_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1775_ _2587_/Q _2584_/Q VGND VGND VPWR VPWR _1777_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2329_/A VGND VGND VPWR VPWR _2327_/Y sky130_fd_sc_hd__inv_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2258_ _2272_/A _2475_/Q VGND VGND VPWR VPWR _2258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ _1608_/B VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2189_ _2231_/A VGND VGND VPWR VPWR _2189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2331__A _2355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2601__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input17_A wbs_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2241__A _2241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1560_ _1560_/A VGND VGND VPWR VPWR _2419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1491_ _2458_/Q _2459_/Q _1495_/S VGND VGND VPWR VPWR _1492_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2112_ _2490_/Q _2111_/X _2078_/X _2101_/X VGND VGND VPWR VPWR _2112_/X sky130_fd_sc_hd__o31a_1
XFILLER_95_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2043_ _2038_/Y _2040_/Y _2042_/X VGND VGND VPWR VPWR _2043_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_48_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1827_ _1722_/X _1828_/C _1828_/D _1828_/B VGND VGND VPWR VPWR _1829_/A sky130_fd_sc_hd__o22a_1
XFILLER_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1758_ _1754_/X _1755_/Y _1789_/C _2437_/Q VGND VGND VPWR VPWR _1759_/B sky130_fd_sc_hd__and4bb_1
XFILLER_102_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1689_ _2415_/Q VGND VGND VPWR VPWR _1693_/C sky130_fd_sc_hd__inv_2
XANTENNA__1990__A _1993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A wbs_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2326__A _2329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2061__A _2083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2236__A _2264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1612_ _2447_/Q _2446_/Q _1612_/C VGND VGND VPWR VPWR _1614_/A sky130_fd_sc_hd__nand3_1
XFILLER_12_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2592_ _2595_/CLK _2592_/D _2357_/Y VGND VGND VPWR VPWR _2592_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_1_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1543_ input44/X _2426_/Q _1545_/S VGND VGND VPWR VPWR _1544_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1474_ _1474_/A VGND VGND VPWR VPWR _2466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1340__A1 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2026_ _2026_/A VGND VGND VPWR VPWR _2294_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1985__A _1987_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1331__A1 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1895__A _1913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1190_ _1324_/A VGND VGND VPWR VPWR _2237_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 wbs_adr_i[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1678__A1_N _1647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2575_ _2577_/CLK _2575_/D _2336_/Y VGND VGND VPWR VPWR _2575_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1526_ input53/X _2434_/Q _1534_/S VGND VGND VPWR VPWR _1527_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1457_ _1457_/A VGND VGND VPWR VPWR _2474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1388_ _1388_/A VGND VGND VPWR VPWR _2505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2009_ _2011_/A VGND VGND VPWR VPWR _2009_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2492__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2360_ _2360_/A VGND VGND VPWR VPWR _2360_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1311_ _1339_/A VGND VGND VPWR VPWR _1311_/X sky130_fd_sc_hd__buf_2
XFILLER_135_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2291_ _2545_/Q VGND VGND VPWR VPWR _2291_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1242_ _1293_/A VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1173_ _1173_/A _1173_/B VGND VGND VPWR VPWR _1177_/A sky130_fd_sc_hd__nor2_2
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2143__B _2236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2558_ _2560_/CLK _2558_/D _2315_/Y VGND VGND VPWR VPWR _2558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1509_ _1509_/A VGND VGND VPWR VPWR _2450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2489_ _2560_/CLK _2489_/D _1984_/Y VGND VGND VPWR VPWR _2489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2262__A2 _2246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2053__B _2061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input47_A wbs_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2228__B _2228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1559__S _1567_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _1863_/A VGND VGND VPWR VPWR _1860_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput12 wbs_adr_i[19] VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1791_ _2591_/Q _2588_/Q _1790_/B VGND VGND VPWR VPWR _2591_/D sky130_fd_sc_hd__a21o_1
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 wbs_adr_i[29] VGND VGND VPWR VPWR _1172_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput34 wbs_cyc_i VGND VGND VPWR VPWR _1165_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 wbs_dat_i[19] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 wbs_dat_i[29] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput67 wbs_stb_i VGND VGND VPWR VPWR _1165_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2412_ _2549_/CLK _2412_/D _1887_/Y VGND VGND VPWR VPWR _2412_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2343_ _2355_/A VGND VGND VPWR VPWR _2348_/A sky130_fd_sc_hd__buf_2
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2274_ _2509_/Q _2241_/X _2252_/X _2032_/X VGND VGND VPWR VPWR _2274_/X sky130_fd_sc_hd__o31a_1
XFILLER_26_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1225_ input54/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__o21ba_1
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1989_ _1993_/A VGND VGND VPWR VPWR _1989_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1993__A _1993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2180__A1 _1621_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2329__A _2329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1233__A _1608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2530__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2064__A _2099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1408__A _1430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2239__A _2272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1912_ _1912_/A VGND VGND VPWR VPWR _1912_/Y sky130_fd_sc_hd__inv_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1843_ _1844_/A VGND VGND VPWR VPWR _1843_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1774_ _2587_/Q _2584_/Q VGND VGND VPWR VPWR _1777_/D sky130_fd_sc_hd__and2_1
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1318__A _1512_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2329_/A VGND VGND VPWR VPWR _2326_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _2257_/A _2292_/B VGND VGND VPWR VPWR _2257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1208_ _1497_/A VGND VGND VPWR VPWR _1608_/B sky130_fd_sc_hd__buf_2
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ _1828_/C _2186_/X _2162_/X _2187_/Y VGND VGND VPWR VPWR _2188_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1988__A _2006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2553__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1898__A _1900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1195__A2 _1191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2426__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1490_ _1490_/A VGND VGND VPWR VPWR _2459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1572__S _1578_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _2241_/A VGND VGND VPWR VPWR _2111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2576__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2042_ _2482_/Q _1346_/A _2016_/X _2246_/A VGND VGND VPWR VPWR _2042_/X sky130_fd_sc_hd__o31a_1
XFILLER_3_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1826_ _2369_/Q _2600_/Q VGND VGND VPWR VPWR _1828_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2151__B _2161_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1757_ _2546_/Q VGND VGND VPWR VPWR _1789_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1688_ _2389_/Q _2386_/Q _1687_/B VGND VGND VPWR VPWR _2389_/D sky130_fd_sc_hd__a21o_1
XFILLER_172_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2311_/A VGND VGND VPWR VPWR _2309_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2449__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2061__B _2061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2599__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2236__B _2236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1567__S _1567_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2252__A _2252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1611_ _2446_/Q _1612_/C _1610_/Y VGND VGND VPWR VPWR _2446_/D sky130_fd_sc_hd__a21oi_1
X_2591_ _2595_/CLK _2591_/D _2356_/Y VGND VGND VPWR VPWR _2591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1542_ _1542_/A VGND VGND VPWR VPWR _2427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1473_ _2466_/Q _2467_/Q _1473_/S VGND VGND VPWR VPWR _1474_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2025_ _2237_/A VGND VGND VPWR VPWR _2292_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2162__A _2249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1809_ _1809_/A _1809_/B VGND VGND VPWR VPWR _2596_/D sky130_fd_sc_hd__nor2_1
XFILLER_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2337__A _2355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2044__B1 _2043_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2072__A _2294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2247__A _2247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2283__B1 _2282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2035__B1 _2034_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2574_ _2576_/CLK _2574_/D _2335_/Y VGND VGND VPWR VPWR _2574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1525_ _1558_/A VGND VGND VPWR VPWR _1534_/S sky130_fd_sc_hd__buf_2
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1456_ _2474_/Q _2475_/Q _1462_/S VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1387_ _2505_/Q _2506_/Q _1395_/S VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2008_ _2011_/A VGND VGND VPWR VPWR _2008_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2274__B1 _2032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1996__A _1999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1236__A _2247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2017__B1 _2513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _2558_/Q _1286_/X _1307_/X _1309_/Y VGND VGND VPWR VPWR _2557_/D sky130_fd_sc_hd__a22o_1
XFILLER_123_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2290_ _2284_/Y _2116_/A _2289_/Y VGND VGND VPWR VPWR _2544_/D sky130_fd_sc_hd__o21ai_2
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ input51/X _1219_/X _1224_/X VGND VGND VPWR VPWR _1241_/X sky130_fd_sc_hd__o21ba_1
XFILLER_61_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1172_ _1172_/A _1172_/B _1172_/C VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__nand3_4
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 _2522_/Q VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_192_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2557_ _2560_/CLK _2557_/D _2314_/Y VGND VGND VPWR VPWR _2557_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1508_ _2450_/Q _2451_/Q _1589_/A VGND VGND VPWR VPWR _1509_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2488_ _2560_/CLK _2488_/D _1983_/Y VGND VGND VPWR VPWR _2488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1439_ _2481_/Q _2482_/Q _1439_/S VGND VGND VPWR VPWR _1440_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1298__A1 input39/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 wbs_adr_i[1] VGND VGND VPWR VPWR _1179_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1790_ _1790_/A _1790_/B VGND VGND VPWR VPWR _2590_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput24 wbs_adr_i[2] VGND VGND VPWR VPWR _1200_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput35 wbs_dat_i[0] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput46 wbs_dat_i[1] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_4
Xinput57 wbs_dat_i[2] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_2
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 wbs_we_i VGND VGND VPWR VPWR _2012_/B sky130_fd_sc_hd__buf_2
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2411_ _2549_/CLK _2411_/D _1886_/Y VGND VGND VPWR VPWR _2411_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2342_ _2342_/A VGND VGND VPWR VPWR _2342_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2273_ _1221_/Y _2237_/X _2249_/X _2272_/Y VGND VGND VPWR VPWR _2273_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_211_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1224_ _1589_/A VGND VGND VPWR VPWR _1224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ _2006_/A VGND VGND VPWR VPWR _1993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2170__A _2170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2482__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2180__A2 _2118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1514__A _1558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2239__B _2473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1911_ _1912_/A VGND VGND VPWR VPWR _1911_/Y sky130_fd_sc_hd__inv_2
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1842_ _1844_/A VGND VGND VPWR VPWR _1842_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1773_ _2434_/Q VGND VGND VPWR VPWR _1777_/C sky130_fd_sc_hd__clkinv_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2329_/A VGND VGND VPWR VPWR _2325_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _2540_/Q VGND VGND VPWR VPWR _2256_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1207_ _1293_/A _2061_/B _1206_/Y VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2187_ _2187_/A _2467_/Q VGND VGND VPWR VPWR _2187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2378__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2075__A _2099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1419__A _1430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _1321_/Y _2062_/X _2074_/X _2109_/Y VGND VGND VPWR VPWR _2110_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2041_ _2146_/A VGND VGND VPWR VPWR _2246_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1825_ _2369_/Q _2600_/Q VGND VGND VPWR VPWR _1828_/D sky130_fd_sc_hd__and2_1
XFILLER_163_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1747_/X _2437_/Q _1754_/X _1755_/Y VGND VGND VPWR VPWR _1759_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1687_ _1687_/A _1687_/B VGND VGND VPWR VPWR _2388_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2520__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2311_/A VGND VGND VPWR VPWR _2308_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1999__A _1999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2239_ _2272_/A _2473_/Q VGND VGND VPWR VPWR _2239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A wbs_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1702__A _1747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1610_ _2446_/Q _1612_/C _1588_/X _1586_/X _1614_/C VGND VGND VPWR VPWR _1610_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_199_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ _2595_/CLK _2590_/D _2354_/Y VGND VGND VPWR VPWR _2590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output90_A _2542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1541_ input45/X _2427_/Q _1545_/S VGND VGND VPWR VPWR _1542_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1583__S _1583_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2543__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1472_ _1472_/A VGND VGND VPWR VPWR _2467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2024_ _2285_/A _2024_/B _2408_/Q VGND VGND VPWR VPWR _2024_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1808_ _1805_/X _1806_/Y _1821_/C _2429_/Q VGND VGND VPWR VPWR _1809_/B sky130_fd_sc_hd__and4bb_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1739_ _1737_/X _2405_/D VGND VGND VPWR VPWR _1740_/A sky130_fd_sc_hd__and2b_1
XFILLER_172_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1493__S _1495_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2416__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2566__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1578__S _1578_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2263__A _2541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2573_ _2576_/CLK _2573_/D _2334_/Y VGND VGND VPWR VPWR _2573_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1524_ _1524_/A VGND VGND VPWR VPWR _2435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1455_ _1455_/A VGND VGND VPWR VPWR _2475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1386_ _1430_/A VGND VGND VPWR VPWR _1395_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2007_ _2011_/A VGND VGND VPWR VPWR _2007_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2589__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1537__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1252__A _1374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2017__A1 _1214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2083__A _2083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1528__A0 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1240_ _2572_/Q _1233_/X _1234_/X _1239_/Y VGND VGND VPWR VPWR _2571_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1171_ _1171_/A _1171_/B VGND VGND VPWR VPWR _1172_/C sky130_fd_sc_hd__nor2_2
XANTENNA__2258__A _2272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1231__A2 _1214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1519__A0 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput101 _2523_/Q VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_192_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2556_ _2560_/CLK _2556_/D _2313_/Y VGND VGND VPWR VPWR _2556_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1507_ _1507_/A VGND VGND VPWR VPWR _2451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2487_ _2549_/CLK _2487_/D _1980_/Y VGND VGND VPWR VPWR _2487_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1438_ _1438_/A VGND VGND VPWR VPWR _2482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1369_ _2547_/Q _1194_/X _1364_/X _1368_/Y VGND VGND VPWR VPWR _2546_/D sky130_fd_sc_hd__a22o_1
XFILLER_210_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1222__A2 _1214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 wbs_adr_i[20] VGND VGND VPWR VPWR _1173_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 wbs_adr_i[30] VGND VGND VPWR VPWR _1171_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput36 wbs_dat_i[10] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput47 wbs_dat_i[20] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput58 wbs_dat_i[30] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2410_ _2553_/CLK _2410_/D _1885_/Y VGND VGND VPWR VPWR _2410_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2341_ _2342_/A VGND VGND VPWR VPWR _2341_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2272_ _2272_/A _2477_/Q VGND VGND VPWR VPWR _2272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1223_ _2575_/Q _1209_/X _1220_/X _1222_/Y VGND VGND VPWR VPWR _2574_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1987_ _1987_/A VGND VGND VPWR VPWR _1987_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2539_ _2569_/CLK _2539_/D VGND VGND VPWR VPWR _2539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2361__A _2361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input52_A wbs_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1910_ _1912_/A VGND VGND VPWR VPWR _1910_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _1844_/A VGND VGND VPWR VPWR _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2271__A _2285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1772_ _2585_/Q _2582_/Q _1771_/B VGND VGND VPWR VPWR _2585_/D sky130_fd_sc_hd__a21o_1
XFILLER_200_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2324_/A VGND VGND VPWR VPWR _2329_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2255_ _2245_/Y _2246_/X _2254_/Y VGND VGND VPWR VPWR _2539_/D sky130_fd_sc_hd__o21ai_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1206_ _2576_/Q VGND VGND VPWR VPWR _1206_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2186_ _2186_/A VGND VGND VPWR VPWR _2186_/X sky130_fd_sc_hd__buf_2
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1350__A _2170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1364__B1_N _1372_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1525__A _1558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2040_ _1361_/Y _2292_/B _2030_/X _2039_/Y VGND VGND VPWR VPWR _2040_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_181_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1170__A _2014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2472__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1824_ _2426_/Q VGND VGND VPWR VPWR _1828_/C sky130_fd_sc_hd__inv_2
XFILLER_34_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1755_ _2581_/Q _2578_/Q VGND VGND VPWR VPWR _1755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1686_ _1777_/A _1686_/B _1686_/C _1686_/D VGND VGND VPWR VPWR _1687_/B sky130_fd_sc_hd__nor4_1
XANTENNA__1591__A1 _1194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2311_/A VGND VGND VPWR VPWR _2307_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2238_ _2238_/A VGND VGND VPWR VPWR _2272_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2169_ _2530_/Q VGND VGND VPWR VPWR _2169_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2498__RESET_B _1995_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1241__B1_N _1224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2495__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A wbs_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2295__C1 _2294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _1540_/A VGND VGND VPWR VPWR _2428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1471_ _2467_/Q _2468_/Q _1473_/S VGND VGND VPWR VPWR _1472_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2023_ _2213_/A VGND VGND VPWR VPWR _2285_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ _1652_/C _2429_/Q _1805_/X _1806_/Y VGND VGND VPWR VPWR _1809_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2368__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1738_ _1821_/C _2439_/Q _2405_/Q VGND VGND VPWR VPWR _2405_/D sky130_fd_sc_hd__a21o_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1669_ _2385_/Q _2382_/Q VGND VGND VPWR VPWR _1673_/D sky130_fd_sc_hd__and2_1
XFILLER_28_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input7_A wbs_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2044__A2 _2022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2283__A2 _2246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2035__A2 _2022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2510__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2572_ _2576_/CLK _2572_/D _2333_/Y VGND VGND VPWR VPWR _2572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1523_ input54/X _2435_/Q _1523_/S VGND VGND VPWR VPWR _1524_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1454_ _2475_/Q _2476_/Q _1462_/S VGND VGND VPWR VPWR _1455_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1385_ _2448_/Q VGND VGND VPWR VPWR _1430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2006_ _2006_/A VGND VGND VPWR VPWR _2011_/A sky130_fd_sc_hd__buf_2
XFILLER_64_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2533__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2017__A2 _2016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2083__B _2134_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1776__A1 _1722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1170_ _2014_/A _1170_/B VGND VGND VPWR VPWR _1512_/A sky130_fd_sc_hd__nor2_4
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1519__A1 _2437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2555_ _2560_/CLK _2555_/D _2311_/Y VGND VGND VPWR VPWR _2555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1506_ _2451_/Q _2452_/Q _1506_/S VGND VGND VPWR VPWR _1507_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2406__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2486_ _2560_/CLK _2486_/D _1979_/Y VGND VGND VPWR VPWR _2486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1437_ _2482_/Q _2483_/Q _1439_/S VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1368_ _1346_/X _2061_/B _1643_/A VGND VGND VPWR VPWR _1368_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2556__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1299_ _2559_/Q VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1263__A _2024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 wbs_adr_i[21] VGND VGND VPWR VPWR _1173_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput26 wbs_adr_i[31] VGND VGND VPWR VPWR _1171_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput37 wbs_dat_i[11] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput48 wbs_dat_i[21] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 wbs_dat_i[31] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_4
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2340_ _2342_/A VGND VGND VPWR VPWR _2340_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2271_ _2285_/A _2285_/B _2436_/Q VGND VGND VPWR VPWR _2271_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_26_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2579__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1222_ _1212_/X _1214_/X _1221_/Y VGND VGND VPWR VPWR _1222_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1901__A _1913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ _1987_/A VGND VGND VPWR VPWR _1986_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2538_ _2569_/CLK _2538_/D VGND VGND VPWR VPWR _2538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2469_ _2595_/CLK _2469_/D _1959_/Y VGND VGND VPWR VPWR _2469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input45_A wbs_dat_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1840_ _1844_/A VGND VGND VPWR VPWR _1840_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2271__B _2285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1771_ _1771_/A _1771_/B VGND VGND VPWR VPWR _2584_/D sky130_fd_sc_hd__nor2_1
XFILLER_204_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2323_/A VGND VGND VPWR VPWR _2323_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2248_/Y _2251_/Y _2253_/X VGND VGND VPWR VPWR _2254_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1205_ _2238_/A VGND VGND VPWR VPWR _2061_/B sky130_fd_sc_hd__buf_2
X_2185_ _2185_/A _2228_/B VGND VGND VPWR VPWR _2185_/Y sky130_fd_sc_hd__nor2_1
XFILLER_187_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1969_ _1975_/A VGND VGND VPWR VPWR _1974_/A sky130_fd_sc_hd__buf_2
XFILLER_33_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2091__B _2161_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ _2601_/Q _2598_/Q _1822_/B VGND VGND VPWR VPWR _2601_/D sky130_fd_sc_hd__a21o_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1754_ _2581_/Q _2578_/Q VGND VGND VPWR VPWR _1754_/X sky130_fd_sc_hd__and2_1
XFILLER_69_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1685_ _1631_/X _1686_/C _1686_/D _1686_/B VGND VGND VPWR VPWR _1687_/A sky130_fd_sc_hd__o22a_1
XANTENNA__1591__A2 _1191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2324_/A VGND VGND VPWR VPWR _2311_/A sky130_fd_sc_hd__buf_2
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2237_ _2237_/A VGND VGND VPWR VPWR _2237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _2159_/Y _2160_/X _2167_/Y VGND VGND VPWR VPWR _2529_/D sky130_fd_sc_hd__o21ai_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2099_ _2099_/A _2457_/Q VGND VGND VPWR VPWR _2099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1536__A _1558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1334__A2 _1311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2295__B1 _2074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1470_ _1470_/A VGND VGND VPWR VPWR _2468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2277__A _2543_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2022_ _2116_/A VGND VGND VPWR VPWR _2022_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2560__RESET_B _2317_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1806_ _2597_/Q _2594_/Q VGND VGND VPWR VPWR _1806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1737_ _1821_/C _2439_/Q _2405_/Q VGND VGND VPWR VPWR _1737_/X sky130_fd_sc_hd__and3_1
XFILLER_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1668_ _2418_/Q VGND VGND VPWR VPWR _1673_/C sky130_fd_sc_hd__inv_2
XFILLER_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1599_ _1599_/A VGND VGND VPWR VPWR _2442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1316__A2 _1311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2462__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2571_ _2576_/CLK _2571_/D _2332_/Y VGND VGND VPWR VPWR _2571_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1522_ _1522_/A VGND VGND VPWR VPWR _2436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1453_ _1486_/A VGND VGND VPWR VPWR _1462_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1384_ _1384_/A VGND VGND VPWR VPWR _2506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2005_ _2005_/A VGND VGND VPWR VPWR _2005_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1234__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2485__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1225__A1 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1776__A2 _1777_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2110__C1 _2109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2554_ _2560_/CLK _2554_/D _2310_/Y VGND VGND VPWR VPWR _2554_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1505_ _1505_/A VGND VGND VPWR VPWR _2452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2485_ _2549_/CLK _2485_/D _1978_/Y VGND VGND VPWR VPWR _2485_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1436_ _1436_/A VGND VGND VPWR VPWR _2483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1367_ _1672_/A VGND VGND VPWR VPWR _1643_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1298_ input39/X _1297_/X _1277_/X VGND VGND VPWR VPWR _1298_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2500__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 wbs_adr_i[22] VGND VGND VPWR VPWR _1174_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 wbs_adr_i[3] VGND VGND VPWR VPWR _2013_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput38 wbs_dat_i[12] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput49 wbs_dat_i[22] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2270_ _2542_/Q VGND VGND VPWR VPWR _2270_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1221_ _2574_/Q VGND VGND VPWR VPWR _1221_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2285__A _2285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1985_ _1987_/A VGND VGND VPWR VPWR _1985_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2537_ _2569_/CLK _2537_/D VGND VGND VPWR VPWR _2537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2523__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2468_ _2601_/CLK _2468_/D _1958_/Y VGND VGND VPWR VPWR _2468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1419_ _1430_/A VGND VGND VPWR VPWR _1428_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2399_ _2459_/CLK _2399_/D _1872_/Y VGND VGND VPWR VPWR _2399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2195__A _2238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input38_A wbs_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ _1767_/X _1768_/Y _1789_/C _2435_/Q VGND VGND VPWR VPWR _1771_/B sky130_fd_sc_hd__and4bb_1
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2546__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _2323_/A VGND VGND VPWR VPWR _2322_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2506_/Q _2241_/X _2252_/X _2231_/X VGND VGND VPWR VPWR _2253_/X sky130_fd_sc_hd__o31a_1
XFILLER_26_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1912__A _1912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1204_ _2026_/A VGND VGND VPWR VPWR _2238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2184_ _2532_/Q VGND VGND VPWR VPWR _2184_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ _1968_/A VGND VGND VPWR VPWR _1968_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1899_ _1900_/A VGND VGND VPWR VPWR _1899_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1594__B1 _1194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1750__A2_N _2438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2419__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2569__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2129__A2 _2062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1718__A2_N _2411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1822_ _1822_/A _1822_/B VGND VGND VPWR VPWR _2600_/D sky130_fd_sc_hd__nor2_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1753_ _2579_/Q _2404_/Q _1752_/B VGND VGND VPWR VPWR _2579_/D sky130_fd_sc_hd__a21o_1
XANTENNA__1576__A0 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1907__A _1913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1684_ _2389_/Q _2386_/Q VGND VGND VPWR VPWR _1686_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2305_/A VGND VGND VPWR VPWR _2305_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2236_ _2264_/A _2236_/B _2432_/Q VGND VGND VPWR VPWR _2236_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_22_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2167_ _2161_/Y _2164_/Y _2166_/X VGND VGND VPWR VPWR _2167_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _2098_/A _2161_/B VGND VGND VPWR VPWR _2098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1567__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1727__A _1777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output69_A _2513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2021_ _2146_/A VGND VGND VPWR VPWR _2116_/A sky130_fd_sc_hd__buf_4
XFILLER_23_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2293__A _2439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1805_ _2597_/Q _2594_/Q VGND VGND VPWR VPWR _1805_/X sky130_fd_sc_hd__and2_1
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ _2546_/Q VGND VGND VPWR VPWR _1821_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1667_ _2383_/Q _2380_/Q _1666_/B VGND VGND VPWR VPWR _2383_/D sky130_fd_sc_hd__a21o_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1598_ _1596_/X _1614_/C _1598_/C VGND VGND VPWR VPWR _1599_/A sky130_fd_sc_hd__and3b_1
XFILLER_63_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2219_ _2212_/Y _2203_/X _2218_/Y VGND VGND VPWR VPWR _2535_/D sky130_fd_sc_hd__o21ai_1
XFILLER_22_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1547__A _1558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1713__C _1751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A wbs_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2570_ _2576_/CLK _2570_/D _2329_/Y VGND VGND VPWR VPWR _2570_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1521_ input55/X _2436_/Q _1523_/S VGND VGND VPWR VPWR _1522_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1452_ _1452_/A VGND VGND VPWR VPWR _2476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1383_ _2506_/Q _2507_/Q _1383_/S VGND VGND VPWR VPWR _1384_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2259__A1 _1777_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2004_ _2005_/A VGND VGND VPWR VPWR _2004_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1719_ _1716_/X _1717_/Y _1751_/C _2411_/Q VGND VGND VPWR VPWR _1720_/B sky130_fd_sc_hd__and4bb_1
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2198__A _2241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1277__A _1374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input68_A wbs_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2110__B1 _2074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1216__A2 _1214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2553_ _2553_/CLK _2553_/D _2309_/Y VGND VGND VPWR VPWR _2553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1504_ _2452_/Q _2453_/Q _1506_/S VGND VGND VPWR VPWR _1505_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2484_ _2560_/CLK _2484_/D _1977_/Y VGND VGND VPWR VPWR _2484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1435_ _2483_/Q _2484_/Q _1439_/S VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1366_ _1722_/A VGND VGND VPWR VPWR _1672_/A sky130_fd_sc_hd__buf_2
XFILLER_112_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1297_ _1297_/A VGND VGND VPWR VPWR _1297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2452__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1207__A2 _2061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput17 wbs_adr_i[23] VGND VGND VPWR VPWR _1174_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput28 wbs_adr_i[4] VGND VGND VPWR VPWR _1167_/B sky130_fd_sc_hd__clkbuf_1
Xinput39 wbs_dat_i[13] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1220_ input55/X _1219_/X _1339_/A VGND VGND VPWR VPWR _1220_/X sky130_fd_sc_hd__o21ba_1
XFILLER_113_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1685__A2 _1686_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2475__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2285__B _2285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1984_ _1987_/A VGND VGND VPWR VPWR _1984_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2536_ _2569_/CLK _2536_/D VGND VGND VPWR VPWR _2536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2467_ _2601_/CLK _2467_/D _1956_/Y VGND VGND VPWR VPWR _2467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418_ _1418_/A VGND VGND VPWR VPWR _2491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2398_ _2459_/CLK _2398_/D _1871_/Y VGND VGND VPWR VPWR _2398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1349_ _2551_/Q _1339_/X _1345_/X _1348_/Y VGND VGND VPWR VPWR _2550_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1364__A1 input35/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2498__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2321_ _2323_/A VGND VGND VPWR VPWR _2321_/Y sky130_fd_sc_hd__inv_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2252_ _2252_/A VGND VGND VPWR VPWR _2252_/X sky130_fd_sc_hd__clkbuf_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1203_ _1512_/A _2028_/B _2028_/C VGND VGND VPWR VPWR _2026_/A sky130_fd_sc_hd__nand3_2
XFILLER_38_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2183_ _2177_/Y _2160_/X _2182_/Y VGND VGND VPWR VPWR _2531_/D sky130_fd_sc_hd__o21ai_1
XFILLER_22_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1967_ _1968_/A VGND VGND VPWR VPWR _1967_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1898_ _1900_/A VGND VGND VPWR VPWR _1898_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2519_ _2553_/CLK _2519_/D VGND VGND VPWR VPWR _2519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input50_A wbs_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2065__A2 _2062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2513__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ _1818_/X _1819_/Y _1821_/C _2427_/Q VGND VGND VPWR VPWR _1822_/B sky130_fd_sc_hd__and4bb_1
XFILLER_34_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1752_ _1752_/A _1752_/B VGND VGND VPWR VPWR _2578_/D sky130_fd_sc_hd__nor2_1
XFILLER_195_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1576__A1 _2411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1683_ _2389_/Q _2386_/Q VGND VGND VPWR VPWR _1686_/D sky130_fd_sc_hd__and2_1
XFILLER_144_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2305_/A VGND VGND VPWR VPWR _2304_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2538_/Q VGND VGND VPWR VPWR _2235_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2166_ _2496_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2166_/X sky130_fd_sc_hd__o31a_1
XFILLER_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2097_ _2522_/Q VGND VGND VPWR VPWR _2097_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2295__A2 _2186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2536__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ _2231_/A VGND VGND VPWR VPWR _2146_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1804_ _2595_/Q _2592_/Q _1803_/B VGND VGND VPWR VPWR _2595_/D sky130_fd_sc_hd__a21o_1
XFILLER_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1735_ _2403_/Q _2400_/Q _1734_/B VGND VGND VPWR VPWR _2403_/D sky130_fd_sc_hd__a21o_1
XFILLER_195_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2409__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1666_ _1666_/A _1666_/B VGND VGND VPWR VPWR _2382_/D sky130_fd_sc_hd__nor2_1
XFILLER_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1597_ _1588_/A _1593_/A _2442_/Q VGND VGND VPWR VPWR _1598_/C sky130_fd_sc_hd__a21o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2559__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2218_ _2214_/Y _2216_/Y _2217_/X VGND VGND VPWR VPWR _2218_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2149_ _2141_/Y _2116_/X _2148_/Y VGND VGND VPWR VPWR _2527_/D sky130_fd_sc_hd__o21ai_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A wbs_adr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1502__S _1506_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1520_ _1520_/A VGND VGND VPWR VPWR _2437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output81_A _2515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1451_ _2476_/Q _2477_/Q _1451_/S VGND VGND VPWR VPWR _1452_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1382_ _1382_/A VGND VGND VPWR VPWR _2507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2259__A2 _2186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2003_ _2005_/A VGND VGND VPWR VPWR _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1718_ _1702_/X _2411_/Q _1716_/X _1717_/Y VGND VGND VPWR VPWR _1720_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1649_ _2379_/Q _2376_/Q VGND VGND VPWR VPWR _1649_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2381__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input5_A wbs_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1458__A0 _2473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1558__A _1558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1449__A0 _2477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2552_ _2560_/CLK _2552_/D _2308_/Y VGND VGND VPWR VPWR _2552_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ _1503_/A VGND VGND VPWR VPWR _2453_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2299__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2483_ _2560_/CLK _2483_/D _1976_/Y VGND VGND VPWR VPWR _2483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1434_ _1434_/A VGND VGND VPWR VPWR _2484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1365_ _2546_/Q VGND VGND VPWR VPWR _1722_/A sky130_fd_sc_hd__inv_2
XFILLER_25_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1296_ _2561_/Q _1286_/X _1292_/X _1295_/Y VGND VGND VPWR VPWR _2560_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2002__A _2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1288__A _2024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1719__C _1751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput18 wbs_adr_i[24] VGND VGND VPWR VPWR _1175_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 wbs_adr_i[5] VGND VGND VPWR VPWR _1167_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_182_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1983_ _1987_/A VGND VGND VPWR VPWR _1983_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1198__A _1497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2535_ _2569_/CLK _2535_/D VGND VGND VPWR VPWR _2535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2466_ _2601_/CLK _2466_/D _1955_/Y VGND VGND VPWR VPWR _2466_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1417_ _2491_/Q _2492_/Q _1417_/S VGND VGND VPWR VPWR _1418_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2397_ _2459_/CLK _2397_/D _1869_/Y VGND VGND VPWR VPWR _2397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1348_ _1346_/X _1341_/X _1347_/Y VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1279_ _2563_/Q VGND VGND VPWR VPWR _2178_/A sky130_fd_sc_hd__inv_2
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1510__S _1589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2323_/A VGND VGND VPWR VPWR _2320_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2442__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _1238_/Y _2237_/X _2249_/X _2250_/Y VGND VGND VPWR VPWR _2251_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_26_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ _2241_/A VGND VGND VPWR VPWR _1293_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2182_ _2178_/Y _2180_/Y _2181_/X VGND VGND VPWR VPWR _2182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2592__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_wb_clk_i clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR _2459_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_181_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1966_ _1968_/A VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2240__B1 _2205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1897_ _1900_/A VGND VGND VPWR VPWR _1897_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2518_ _2553_/CLK _2518_/D VGND VGND VPWR VPWR _2518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2449_ _2549_/CLK _2449_/D _1934_/Y VGND VGND VPWR VPWR _2449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1282__A1 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2465__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A wbs_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1820_ _1652_/C _2427_/Q _1818_/X _1819_/Y VGND VGND VPWR VPWR _1822_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1751_ _1748_/X _1749_/Y _1751_/C _2438_/Q VGND VGND VPWR VPWR _1752_/B sky130_fd_sc_hd__and4bb_1
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1682_ _2416_/Q VGND VGND VPWR VPWR _1686_/C sky130_fd_sc_hd__inv_2
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2305_/A VGND VGND VPWR VPWR _2303_/Y sky130_fd_sc_hd__inv_2
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2227_/Y _2203_/X _2233_/Y VGND VGND VPWR VPWR _2537_/D sky130_fd_sc_hd__o21ai_1
XFILLER_41_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2165_ _2165_/A VGND VGND VPWR VPWR _2165_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2096_ _2089_/Y _2071_/X _2095_/Y VGND VGND VPWR VPWR _2521_/D sky130_fd_sc_hd__o21ai_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2488__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1949_ _1949_/A VGND VGND VPWR VPWR _1949_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1386__A _1430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2010__A _2011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1727__C _1727_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1803_ _1803_/A _1803_/B VGND VGND VPWR VPWR _2594_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1734_ _1734_/A _1734_/B VGND VGND VPWR VPWR _2402_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1665_ _1662_/X _1663_/Y _1706_/C _2419_/Q VGND VGND VPWR VPWR _1666_/B sky130_fd_sc_hd__and4bb_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1596_ _2441_/Q _2440_/Q _2442_/Q VGND VGND VPWR VPWR _1596_/X sky130_fd_sc_hd__and3_1
XFILLER_193_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2217_ _2502_/Q _2198_/X _2208_/X _2189_/X VGND VGND VPWR VPWR _2217_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2148_ _2143_/Y _2145_/Y _2147_/X VGND VGND VPWR VPWR _2148_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2079_ _2486_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2079_/X sky130_fd_sc_hd__o31a_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2005__A _2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2503__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ _1450_/A VGND VGND VPWR VPWR _2477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output74_A _2527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1381_ _2507_/Q _2508_/Q _1383_/S VGND VGND VPWR VPWR _1382_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2002_ _2005_/A VGND VGND VPWR VPWR _2002_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1467__A1 _2470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1717_ _2399_/Q _2396_/Q VGND VGND VPWR VPWR _1717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2526__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1648_ _2379_/Q _2376_/Q VGND VGND VPWR VPWR _1648_/X sky130_fd_sc_hd__and2_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1579_ _1579_/A VGND VGND VPWR VPWR _2410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1449__A1 _2478_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2110__A2 _2062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1763__A2_N _2436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2549__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1187__C _1187_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2551_ _2553_/CLK _2551_/D _2307_/Y VGND VGND VPWR VPWR _2551_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1502_ _2453_/Q _2454_/Q _1506_/S VGND VGND VPWR VPWR _1503_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2482_ _2512_/CLK _2482_/D _1974_/Y VGND VGND VPWR VPWR _2482_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _2484_/Q _2485_/Q _1439_/S VGND VGND VPWR VPWR _1434_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1364_ input35/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1364_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1295_ _1293_/X _1288_/X _2151_/A VGND VGND VPWR VPWR _1295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1569__A _2186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1719__D _2411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput19 wbs_adr_i[25] VGND VGND VPWR VPWR _1175_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1508__S _1589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2371__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1982_ _2006_/A VGND VGND VPWR VPWR _1987_/A sky130_fd_sc_hd__buf_2
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2534_ _2569_/CLK _2534_/D VGND VGND VPWR VPWR _2534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2465_ _2601_/CLK _2465_/D _1954_/Y VGND VGND VPWR VPWR _2465_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1416_ _1416_/A VGND VGND VPWR VPWR _2492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2396_ _2459_/CLK _2396_/D _1868_/Y VGND VGND VPWR VPWR _2396_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1347_ _2550_/Q VGND VGND VPWR VPWR _1347_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1530__A0 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1278_ input43/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1278_/X sky130_fd_sc_hd__o21ba_1
XFILLER_186_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2013__A _2013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1521__A0 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__C_N _2409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2272_/A _2474_/Q VGND VGND VPWR VPWR _2250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1201_ _1512_/D VGND VGND VPWR VPWR _2241_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2181_ _2498_/Q _2155_/X _2165_/X _2146_/X VGND VGND VPWR VPWR _2181_/X sky130_fd_sc_hd__o31a_1
XFILLER_22_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1965_ _1968_/A VGND VGND VPWR VPWR _1965_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1896_ _1900_/A VGND VGND VPWR VPWR _1896_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2517_ _2553_/CLK _2517_/D VGND VGND VPWR VPWR _2517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2448_ _2549_/CLK _2448_/D _1933_/Y VGND VGND VPWR VPWR _2448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2379_ _2601_/CLK _2379_/D _1847_/Y VGND VGND VPWR VPWR _2379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2008__A _2011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input36_A wbs_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1757__A _2546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1360__B1_N _1372_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1750_ _1747_/X _2438_/Q _1748_/X _1749_/Y VGND VGND VPWR VPWR _1752_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1681_ _2387_/Q _2384_/Q _1680_/B VGND VGND VPWR VPWR _2387_/D sky130_fd_sc_hd__a21o_1
XFILLER_176_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2302_ _2305_/A VGND VGND VPWR VPWR _2302_/Y sky130_fd_sc_hd__inv_2
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2233_ _2228_/Y _2230_/Y _2232_/X VGND VGND VPWR VPWR _2233_/Y sky130_fd_sc_hd__o21ai_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2164_ _1636_/C _2118_/X _2162_/X _2163_/Y VGND VGND VPWR VPWR _2164_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1431__S _1439_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2095_ _2091_/Y _2093_/Y _2094_/X VGND VGND VPWR VPWR _2095_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1948_ _1949_/A VGND VGND VPWR VPWR _1948_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1879_ _1881_/A VGND VGND VPWR VPWR _1879_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2582__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1802_ _1799_/X _1800_/Y _1821_/C _2430_/Q VGND VGND VPWR VPWR _1803_/B sky130_fd_sc_hd__and4bb_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1733_ _1730_/X _1731_/Y _1751_/C _2409_/Q VGND VGND VPWR VPWR _1734_/B sky130_fd_sc_hd__and4bb_1
XFILLER_184_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1664_ _1647_/X _2419_/Q _1662_/X _1663_/Y VGND VGND VPWR VPWR _1666_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1595_ _1588_/A _1593_/A _1594_/Y VGND VGND VPWR VPWR _2441_/D sky130_fd_sc_hd__a21oi_1
XFILLER_8_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2111__A _2241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1950__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2216_ _1258_/Y _2135_/X _2205_/X _2215_/Y VGND VGND VPWR VPWR _2216_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2147_ _2494_/Q _2111_/X _2122_/X _2146_/X VGND VGND VPWR VPWR _2147_/X sky130_fd_sc_hd__o31a_1
XFILLER_167_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2078_ _2165_/A VGND VGND VPWR VPWR _2078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1397__A _1430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1828__C _1828_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1380_ _1380_/A VGND VGND VPWR VPWR _2508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_1_0_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2478__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2001_ _2005_/A VGND VGND VPWR VPWR _2001_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2106__A _2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1716_ _2399_/Q _2396_/Q VGND VGND VPWR VPWR _1716_/X sky130_fd_sc_hd__and2_1
XFILLER_69_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1647_ _1747_/A VGND VGND VPWR VPWR _1647_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ input57/X _2410_/Q _1578_/S VGND VGND VPWR VPWR _1579_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2016__A _2252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ _2553_/CLK _2550_/D _2305_/Y VGND VGND VPWR VPWR _2550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1501_ _1501_/A VGND VGND VPWR VPWR _2454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2481_ _2512_/CLK _2481_/D _1973_/Y VGND VGND VPWR VPWR _2481_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1432_ _1432_/A VGND VGND VPWR VPWR _2485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1363_ _2548_/Q _1339_/X _1360_/X _1362_/Y VGND VGND VPWR VPWR _2547_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ _2560_/Q VGND VGND VPWR VPWR _2151_/A sky130_fd_sc_hd__inv_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input66_A wbs_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1751__C _1751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2516__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1981_ input1/X VGND VGND VPWR VPWR _2006_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ _2569_/CLK _2533_/D VGND VGND VPWR VPWR _2533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2464_ _2601_/CLK _2464_/D _1953_/Y VGND VGND VPWR VPWR _2464_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1415_ _2492_/Q _2493_/Q _1417_/S VGND VGND VPWR VPWR _1416_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2395_ _2459_/CLK _2395_/D _1867_/Y VGND VGND VPWR VPWR _2395_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1346_ _1346_/A VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ _1374_/A VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2086__A2 _2066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1521__A1 _2436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2539__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1200_ _1200_/A VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__inv_2
XFILLER_61_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2180_ _1621_/C _2118_/X _2162_/X _2179_/Y VGND VGND VPWR VPWR _2180_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_211_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1964_ _1968_/A VGND VGND VPWR VPWR _1964_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1895_ _1913_/A VGND VGND VPWR VPWR _1900_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2516_ _2553_/CLK _2516_/D VGND VGND VPWR VPWR _2516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2447_ _2599_/CLK _2447_/D _1931_/Y VGND VGND VPWR VPWR _2447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2378_ _2601_/CLK _2378_/D _1846_/Y VGND VGND VPWR VPWR _2378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1329_ _2555_/Q _1311_/X _1326_/X _1328_/Y VGND VGND VPWR VPWR _2554_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2059__A2 _2022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2216__C1 _2215_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2024__A _2285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2298__A2 _2116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input29_A wbs_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _1680_/A _1680_/B VGND VGND VPWR VPWR _2386_/D sky130_fd_sc_hd__nor2_1
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2301_ _2305_/A VGND VGND VPWR VPWR _2301_/Y sky130_fd_sc_hd__inv_2
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _2504_/Q _2198_/X _2208_/X _2231_/X VGND VGND VPWR VPWR _2232_/X sky130_fd_sc_hd__o31a_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2163_ _2187_/A _2464_/Q VGND VGND VPWR VPWR _2163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2094_ _2488_/Q _2066_/X _2078_/X _2056_/X VGND VGND VPWR VPWR _2094_/X sky130_fd_sc_hd__o31a_1
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2109__A _2144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1947_ _1949_/A VGND VGND VPWR VPWR _1947_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1878_ _1881_/A VGND VGND VPWR VPWR _1878_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2384__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2019__A _2026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ _1652_/C _2430_/Q _1799_/X _1800_/Y VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_34_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _1702_/X _2409_/Q _1730_/X _1731_/Y VGND VGND VPWR VPWR _1734_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_195_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1663_ _2383_/Q _2380_/Q VGND VGND VPWR VPWR _1663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1594_ _1588_/A _1593_/A _1194_/X VGND VGND VPWR VPWR _1594_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2215_ _2229_/A _2470_/Q VGND VGND VPWR VPWR _2215_/Y sky130_fd_sc_hd__nand2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2146_ _2146_/A VGND VGND VPWR VPWR _2146_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2077_ _2252_/A VGND VGND VPWR VPWR _2165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2302__A _2305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2000_ _2006_/A VGND VGND VPWR VPWR _2005_/A sky130_fd_sc_hd__buf_2
XFILLER_23_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1715_ _2397_/Q _2394_/Q _1714_/B VGND VGND VPWR VPWR _2397_/D sky130_fd_sc_hd__a21o_1
XANTENNA__1437__S _1439_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1646_ _2546_/Q VGND VGND VPWR VPWR _1747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1577_ _1577_/A VGND VGND VPWR VPWR _2411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2422__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2572__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2129_ _1308_/Y _2062_/X _2119_/X _2128_/Y VGND VGND VPWR VPWR _2129_/Y sky130_fd_sc_hd__o211ai_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1201__A _1512_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2032__A _2231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input11_A wbs_adr_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1500_ _2454_/Q _2455_/Q _1506_/S VGND VGND VPWR VPWR _1501_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2480_ _2512_/CLK _2480_/D _1972_/Y VGND VGND VPWR VPWR _2480_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2445__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1431_ _2485_/Q _2486_/Q _1439_/S VGND VGND VPWR VPWR _1432_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1362_ _1346_/X _1341_/X _1361_/Y VGND VGND VPWR VPWR _1362_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput90 _2542_/Q VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2595__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1293_ _1293_/A VGND VGND VPWR VPWR _1293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1629_ _1629_/A _1629_/B VGND VGND VPWR VPWR _2372_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input3_A wbs_adr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2027__A _2294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2468__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input59_A wbs_dat_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1751__D _2438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ _1980_/A VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__inv_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2601_ _2601_/CLK _2601_/D _2367_/Y VGND VGND VPWR VPWR _2601_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2532_ _2569_/CLK _2532_/D VGND VGND VPWR VPWR _2532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2463_ _2601_/CLK _2463_/D _1952_/Y VGND VGND VPWR VPWR _2463_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1414_ _1414_/A VGND VGND VPWR VPWR _2493_/D sky130_fd_sc_hd__clkbuf_1
X_2394_ _2459_/CLK _2394_/D _1866_/Y VGND VGND VPWR VPWR _2394_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1345_ input61/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1345_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1276_ _2565_/Q _1261_/X _1273_/X _1275_/Y VGND VGND VPWR VPWR _2564_/D sky130_fd_sc_hd__a22o_1
XFILLER_186_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2086__A3 _2078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1686__A _1777_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1349__A2 _1339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2204__B _2228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1963_ _1975_/A VGND VGND VPWR VPWR _1968_/A sky130_fd_sc_hd__buf_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1894_ _1894_/A VGND VGND VPWR VPWR _1894_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2515_ _2553_/CLK _2515_/D VGND VGND VPWR VPWR _2515_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2446_ _2599_/CLK _2446_/D _1930_/Y VGND VGND VPWR VPWR _2446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2377_ _2601_/CLK _2377_/D _1844_/Y VGND VGND VPWR VPWR _2377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1328_ _1320_/X _1313_/X _2098_/A VGND VGND VPWR VPWR _1328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1259_ _1242_/X _1237_/X _1258_/Y VGND VGND VPWR VPWR _1259_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2216__B1 _2205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2305__A _2305_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2024__B _2024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2506__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2207__B1 _2205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2215__A _2229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ _2324_/A VGND VGND VPWR VPWR _2305_/A sky130_fd_sc_hd__buf_2
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2231_ _2231_/A VGND VGND VPWR VPWR _2231_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2162_ _2249_/A VGND VGND VPWR VPWR _2162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2093_ _1693_/C _1583_/S _2074_/X _2092_/Y VGND VGND VPWR VPWR _2093_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_78_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1946_ _1949_/A VGND VGND VPWR VPWR _1946_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1877_ _1881_/A VGND VGND VPWR VPWR _1877_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2529__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2429_ _2577_/CLK _2429_/D _1909_/Y VGND VGND VPWR VPWR _2429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1204__A _2026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2019__B _2252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1800_ _2595_/Q _2592_/Q VGND VGND VPWR VPWR _1800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1731_ _2403_/Q _2400_/Q VGND VGND VPWR VPWR _1731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1662_ _2383_/Q _2380_/Q VGND VGND VPWR VPWR _1662_/X sky130_fd_sc_hd__and2_1
XFILLER_201_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1593_ _1593_/A _1593_/B VGND VGND VPWR VPWR _2440_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2214_ _2264_/A _2236_/B _2429_/Q VGND VGND VPWR VPWR _2214_/Y sky130_fd_sc_hd__nor3b_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2145_ _1299_/Y _2135_/X _2119_/X _2144_/Y VGND VGND VPWR VPWR _2145_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__1807__A1_N _1652_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2076_ _1342_/Y _2062_/X _2074_/X _2075_/Y VGND VGND VPWR VPWR _2076_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_208_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1929_ _1931_/A VGND VGND VPWR VPWR _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2374__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1714_ _1714_/A _1714_/B VGND VGND VPWR VPWR _2396_/D sky130_fd_sc_hd__nor2_1
XFILLER_195_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1645_ _2377_/Q _2374_/Q _1644_/B VGND VGND VPWR VPWR _2377_/D sky130_fd_sc_hd__a21o_1
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1576_ input60/X _2411_/Q _1578_/S VGND VGND VPWR VPWR _1577_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2104__A2 _2071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _2144_/A _2460_/Q VGND VGND VPWR VPWR _2128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _2052_/Y _2022_/X _2058_/Y VGND VGND VPWR VPWR _2517_/D sky130_fd_sc_hd__o21ai_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2313__A _2317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A VGND VGND VPWR VPWR _1439_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1361_ _2547_/Q VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput80 _2533_/Q VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput91 _2543_/Q VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_190_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1292_ input40/X _1272_/X _1277_/X VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__o21ba_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1302__A _1374_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2117__B _2161_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2595_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1628_ _1643_/A _1628_/B _1628_/C _1628_/D VGND VGND VPWR VPWR _1629_/B sky130_fd_sc_hd__nor4_1
XFILLER_28_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1559_ input37/X _2419_/Q _1567_/S VGND VGND VPWR VPWR _1560_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1827__A1 _1722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2412__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2600_ _2601_/CLK _2600_/D _2366_/Y VGND VGND VPWR VPWR _2600_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2531_ _2569_/CLK _2531_/D VGND VGND VPWR VPWR _2531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2562__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2462_ _2601_/CLK _2462_/D _1949_/Y VGND VGND VPWR VPWR _2462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1413_ _2493_/Q _2494_/Q _1417_/S VGND VGND VPWR VPWR _1414_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1515__A0 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2393_ _2459_/CLK _2393_/D _1865_/Y VGND VGND VPWR VPWR _2393_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1344_ _2552_/Q _1339_/X _1340_/X _1343_/Y VGND VGND VPWR VPWR _2551_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1275_ _1268_/X _1263_/X _2185_/A VGND VGND VPWR VPWR _1275_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2128__A _2144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1506__A0 _2451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2038__A _2083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1877__A _1881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2585__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ _1962_/A VGND VGND VPWR VPWR _1962_/Y sky130_fd_sc_hd__inv_2
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1893_ _1894_/A VGND VGND VPWR VPWR _1893_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2514_ _2553_/CLK _2514_/D VGND VGND VPWR VPWR _2514_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2445_ _2599_/CLK _2445_/D _1929_/Y VGND VGND VPWR VPWR _2445_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2376_ _2601_/CLK _2376_/D _1843_/Y VGND VGND VPWR VPWR _2376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1327_ _2554_/Q VGND VGND VPWR VPWR _2098_/A sky130_fd_sc_hd__inv_2
XFILLER_22_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1258_ _2567_/Q VGND VGND VPWR VPWR _1258_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1189_ _2213_/A _1512_/A _2028_/B _2028_/C VGND VGND VPWR VPWR _1324_/A sky130_fd_sc_hd__nand4_1
XFILLER_129_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2321__A _2323_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2207__A1 _1815_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2215__B _2470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2231__A _2231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _1796_/C _2186_/X _2205_/X _2229_/Y VGND VGND VPWR VPWR _2230_/Y sky130_fd_sc_hd__o211ai_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2600__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2161_ _2161_/A _2161_/B VGND VGND VPWR VPWR _2161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2092_ _2099_/A _2456_/Q VGND VGND VPWR VPWR _2092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1945_ _1949_/A VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1876_ _1882_/A VGND VGND VPWR VPWR _1881_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2141__A _2527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1980__A _1980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2428_ _2576_/CLK _2428_/D _1908_/Y VGND VGND VPWR VPWR _2428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2359_ _2360_/A VGND VGND VPWR VPWR _2359_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2316__A _2317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1890__A _1894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input34_A wbs_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1730_ _2403_/Q _2400_/Q VGND VGND VPWR VPWR _1730_/X sky130_fd_sc_hd__and2_1
XFILLER_157_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1661_ _2381_/Q _2378_/Q _1660_/B VGND VGND VPWR VPWR _2381_/D sky130_fd_sc_hd__a21o_1
XFILLER_176_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1592_ _2440_/Q VGND VGND VPWR VPWR _1593_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2213_/A VGND VGND VPWR VPWR _2264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2144_ _2144_/A _2462_/Q VGND VGND VPWR VPWR _2144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2075_ _2099_/A _2454_/Q VGND VGND VPWR VPWR _2075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2136__A _2144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1975__A _1975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1928_ _1931_/A VGND VGND VPWR VPWR _1928_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ _1863_/A VGND VGND VPWR VPWR _1859_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1770__D _2435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2519__CLK _2553_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1713_ _1709_/X _1710_/Y _1751_/C _2412_/Q VGND VGND VPWR VPWR _1714_/B sky130_fd_sc_hd__and4bb_1
XFILLER_121_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1644_ _1644_/A _1644_/B VGND VGND VPWR VPWR _2376_/D sky130_fd_sc_hd__nor2_1
XFILLER_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1575_ _1575_/A VGND VGND VPWR VPWR _2412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2127_ _2194_/A _2134_/B _2419_/Q VGND VGND VPWR VPWR _2127_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_148_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2058_ _2053_/Y _2055_/Y _2057_/X VGND VGND VPWR VPWR _2058_/Y sky130_fd_sc_hd__o21ai_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2040__A2 _2292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1303__A1 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2031__A2 _2292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1360_ input46/X _2046_/B _1372_/S VGND VGND VPWR VPWR _1360_/X sky130_fd_sc_hd__o21ba_1
Xoutput70 _2514_/Q VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput81 _2515_/Q VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput92 _2516_/Q VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1291_ _2562_/Q _1286_/X _1287_/X _1290_/Y VGND VGND VPWR VPWR _2561_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2491__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1627_ _1828_/A _1628_/C _1628_/D _1628_/B VGND VGND VPWR VPWR _1629_/A sky130_fd_sc_hd__o22a_1
XFILLER_99_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1558_ _1558_/A VGND VGND VPWR VPWR _1567_/S sky130_fd_sc_hd__buf_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1489_ _2459_/Q _2460_/Q _1495_/S VGND VGND VPWR VPWR _1490_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2285__C_N _2438_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2324__A _2324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1827__A2 _1828_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2530_ _2569_/CLK _2530_/D VGND VGND VPWR VPWR _2530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2461_ _2549_/CLK _2461_/D _1948_/Y VGND VGND VPWR VPWR _2461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1412_ _1412_/A VGND VGND VPWR VPWR _2494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2392_ _2459_/CLK _2392_/D _1863_/Y VGND VGND VPWR VPWR _2392_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1515__A1 _2439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1343_ _1320_/X _1341_/X _1342_/Y VGND VGND VPWR VPWR _1343_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1274_ _2564_/Q VGND VGND VPWR VPWR _2185_/A sky130_fd_sc_hd__inv_2
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1313__A _2024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1686__C _1686_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2144__A _2144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1983__A _1987_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1506__A1 _2452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2319__A _2323_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2038__B _2061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2054__A _2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1893__A _1894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input64_A wbs_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2229__A _2229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ _1962_/A VGND VGND VPWR VPWR _1961_/Y sky130_fd_sc_hd__inv_2
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1892_ _1894_/A VGND VGND VPWR VPWR _1892_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2513_ _2553_/CLK _2513_/D VGND VGND VPWR VPWR _2513_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_192_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2444_ _2599_/CLK _2444_/D _1928_/Y VGND VGND VPWR VPWR _2444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2375_ _2601_/CLK _2375_/D _1842_/Y VGND VGND VPWR VPWR _2375_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ input65/X _1325_/X _1302_/X VGND VGND VPWR VPWR _1326_/X sky130_fd_sc_hd__o21ba_1
XFILLER_211_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1257_ input48/X _1246_/X _1252_/X VGND VGND VPWR VPWR _1257_/X sky130_fd_sc_hd__o21ba_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1188_ _1188_/A _1188_/B VGND VGND VPWR VPWR _2028_/C sky130_fd_sc_hd__nor2_4
XFILLER_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1978__A _1980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2216__A2 _2135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1218__A _2237_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1888__A _2361_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2552__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2207__A2 _2186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2160_ _2246_/A VGND VGND VPWR VPWR _2160_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2091_ _2091_/A _2161_/B VGND VGND VPWR VPWR _2091_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1944_ _1944_/A VGND VGND VPWR VPWR _1949_/A sky130_fd_sc_hd__buf_2
XFILLER_202_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1875_ _1875_/A VGND VGND VPWR VPWR _1875_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2425__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2427_ _2576_/CLK _2427_/D _1906_/Y VGND VGND VPWR VPWR _2427_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_170_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2358_ _2360_/A VGND VGND VPWR VPWR _2358_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ _1293_/X _1288_/X _1308_/Y VGND VGND VPWR VPWR _1309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2289_ _2285_/Y _2287_/Y _2288_/X VGND VGND VPWR VPWR _2289_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_61_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A wbs_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1660_ _1660_/A _1660_/B VGND VGND VPWR VPWR _2380_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2448__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1591_ _1194_/X _1191_/X _1593_/B VGND VGND VPWR VPWR _2448_/D sky130_fd_sc_hd__o21ai_1
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2598__CLK _2599_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2535_/Q VGND VGND VPWR VPWR _2212_/Y sky130_fd_sc_hd__inv_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2143_ _2194_/A _2236_/B _2421_/Q VGND VGND VPWR VPWR _2143_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_113_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2074_ _2074_/A VGND VGND VPWR VPWR _2074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ _1931_/A VGND VGND VPWR VPWR _1927_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2152__A _2238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1858_ _1882_/A VGND VGND VPWR VPWR _1863_/A sky130_fd_sc_hd__buf_2
XFILLER_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1789_ _1786_/X _1787_/Y _1789_/C _2432_/Q VGND VGND VPWR VPWR _1790_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__1991__A _1993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2327__A _2329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2062__A _2170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2237__A _2237_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1712_ _1747_/A VGND VGND VPWR VPWR _1751_/C sky130_fd_sc_hd__buf_2
XFILLER_195_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1643_ _1643_/A _1643_/B _1643_/C _1643_/D VGND VGND VPWR VPWR _1644_/B sky130_fd_sc_hd__nor4_1
XFILLER_12_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ input61/X _2412_/Q _1578_/S VGND VGND VPWR VPWR _1575_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2126_ _2525_/Q VGND VGND VPWR VPWR _2126_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2057_ _2484_/Q _1346_/A _2016_/X _2056_/X VGND VGND VPWR VPWR _2057_/X sky130_fd_sc_hd__o31a_1
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1986__A _1987_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1896__A _1900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput71 _2524_/Q VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_29_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput82 _2534_/Q VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput93 _2544_/Q VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_110_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ _1268_/X _1288_/X _2161_/A VGND VGND VPWR VPWR _1290_/Y sky130_fd_sc_hd__o21ai_1
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1570__S _1578_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1626_ _2373_/Q _2370_/Q VGND VGND VPWR VPWR _1628_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1557_ _1557_/A VGND VGND VPWR VPWR _2420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1488_ _1488_/A VGND VGND VPWR VPWR _2460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2109_ _2144_/A _2458_/Q VGND VGND VPWR VPWR _2109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2509__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1460__A1 _2473_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1565__S _1567_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2250__A _2272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2460_ _2601_/CLK _2460_/D _1947_/Y VGND VGND VPWR VPWR _2460_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1411_ _2494_/Q _2495_/Q _1417_/S VGND VGND VPWR VPWR _1412_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2391_ _2459_/CLK _2391_/D _1862_/Y VGND VGND VPWR VPWR _2391_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1342_ _2551_/Q VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1273_ input44/X _1272_/X _1252_/X VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__o21ba_1
XFILLER_81_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1451__A1 _2477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2160__A _2246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1609_ _1609_/A VGND VGND VPWR VPWR _2445_/D sky130_fd_sc_hd__clkbuf_1
X_2589_ _2595_/CLK _2589_/D _2353_/Y VGND VGND VPWR VPWR _2589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input1_A wb_rst_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2054__B _2452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2481__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A wbs_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ _1962_/A VGND VGND VPWR VPWR _1960_/Y sky130_fd_sc_hd__inv_2
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1891_ _1894_/A VGND VGND VPWR VPWR _1891_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2512_ _2512_/CLK _2512_/D _2011_/Y VGND VGND VPWR VPWR _2512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2443_ _2599_/CLK _2443_/D _1927_/Y VGND VGND VPWR VPWR _2443_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2374_ _2601_/CLK _2374_/D _1841_/Y VGND VGND VPWR VPWR _2374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1325_ _2170_/A VGND VGND VPWR VPWR _1325_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1256_ _2569_/Q _1233_/X _1253_/X _1255_/Y VGND VGND VPWR VPWR _2568_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1187_ _1187_/A _1187_/B _1187_/C _1187_/D VGND VGND VPWR VPWR _1188_/B sky130_fd_sc_hd__nand4_4
XFILLER_129_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2155__A _2241_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1994__A _2006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2090_ _2170_/A VGND VGND VPWR VPWR _2161_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2377__CLK _2601_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1943_ _1943_/A VGND VGND VPWR VPWR _1943_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ _1875_/A VGND VGND VPWR VPWR _1874_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1319__A _2066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2426_ _2576_/CLK _2426_/D _1905_/Y VGND VGND VPWR VPWR _2426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2357_ _2360_/A VGND VGND VPWR VPWR _2357_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1308_ _2557_/Q VGND VGND VPWR VPWR _1308_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2288_ _2511_/Q _2066_/A _2165_/A _2032_/X VGND VGND VPWR VPWR _2288_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1989__A _1993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1239_ _1212_/X _1237_/X _1238_/Y VGND VGND VPWR VPWR _1239_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1581__A0 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1899__A _1900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1698__A1_N _1647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1590_ _1586_/X _1588_/X _1614_/C VGND VGND VPWR VPWR _1593_/B sky130_fd_sc_hd__o21ai_1
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output88_A _2540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1572__A0 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2202_/Y _2203_/X _2210_/Y VGND VGND VPWR VPWR _2534_/D sky130_fd_sc_hd__o21ai_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2142_ _2247_/A VGND VGND VPWR VPWR _2236_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2073_ _2083_/A _2134_/B _2413_/Q VGND VGND VPWR VPWR _2073_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1926_ _1944_/A VGND VGND VPWR VPWR _1931_/A sky130_fd_sc_hd__buf_2
XFILLER_202_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1857_ _2361_/A VGND VGND VPWR VPWR _1882_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1788_ _1652_/C _2432_/Q _1786_/X _1787_/Y VGND VGND VPWR VPWR _1790_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2542__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2409_ _2549_/CLK _2409_/D _1884_/Y VGND VGND VPWR VPWR _2409_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1512__A _1512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2343__A _2355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1554__A0 input39/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2415__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1711_ _1702_/X _2412_/Q _1709_/X _1710_/Y VGND VGND VPWR VPWR _1714_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2565__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1642_ _1631_/X _1643_/C _1643_/D _1643_/B VGND VGND VPWR VPWR _1644_/A sky130_fd_sc_hd__o22a_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1573_ _1573_/A VGND VGND VPWR VPWR _2413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2125_ _2115_/Y _2116_/X _2124_/Y VGND VGND VPWR VPWR _2524_/D sky130_fd_sc_hd__o21ai_1
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2056_ _2146_/A VGND VGND VPWR VPWR _2056_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1909_ _1912_/A VGND VGND VPWR VPWR _1909_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2588__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2073__A _2083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput72 _2525_/Q VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput83 _2535_/Q VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 _2545_/Q VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2248__A _2264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1625_ _2373_/Q _2370_/Q VGND VGND VPWR VPWR _1628_/D sky130_fd_sc_hd__and2_1
XFILLER_138_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1556_ input38/X _2420_/Q _1556_/S VGND VGND VPWR VPWR _1557_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1487_ _2460_/Q _2461_/Q _1495_/S VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2108_ _2247_/A VGND VGND VPWR VPWR _2144_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1997__A _1999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2039_ _2054_/A _2450_/Q VGND VGND VPWR VPWR _2039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1237__A _2024_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1410_ _1410_/A VGND VGND VPWR VPWR _2495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2390_ _2459_/CLK _2390_/D _1861_/Y VGND VGND VPWR VPWR _2390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output70_A _2514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1341_ _2054_/A VGND VGND VPWR VPWR _1341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1581__S _1583_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1272_ _1297_/A VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1608_ _1612_/C _1608_/B _1608_/C VGND VGND VPWR VPWR _1609_/A sky130_fd_sc_hd__and3b_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2588_ _2595_/CLK _2588_/D _2352_/Y VGND VGND VPWR VPWR _2588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1539_ input47/X _2428_/Q _1545_/S VGND VGND VPWR VPWR _1540_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1491__S _1495_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1430__A _1430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1890_ _1894_/A VGND VGND VPWR VPWR _1890_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1576__S _1578_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2511_ _2512_/CLK _2511_/D _2010_/Y VGND VGND VPWR VPWR _2511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2442_ _2599_/CLK _2442_/D _1925_/Y VGND VGND VPWR VPWR _2442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2373_ _2601_/CLK _2373_/D _1840_/Y VGND VGND VPWR VPWR _2373_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1324_ _1324_/A VGND VGND VPWR VPWR _2170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1255_ _1242_/X _1237_/X _1254_/Y VGND VGND VPWR VPWR _1255_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_204_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1186_ input8/X input7/X VGND VGND VPWR VPWR _1187_/D sky130_fd_sc_hd__nor2_2
XFILLER_20_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2171__A _2171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1360__A1 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1351__A1 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2256__A _2540_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ _1943_/A VGND VGND VPWR VPWR _1942_/Y sky130_fd_sc_hd__inv_2
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1873_ _1875_/A VGND VGND VPWR VPWR _1873_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2425_ _2576_/CLK _2425_/D _1904_/Y VGND VGND VPWR VPWR _2425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2356_ _2360_/A VGND VGND VPWR VPWR _2356_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1307_ input37/X _1297_/X _1302_/X VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__o21ba_1
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2287_ _1206_/Y _1297_/A _2074_/A _2286_/Y VGND VGND VPWR VPWR _2287_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_61_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1238_ _2571_/Q VGND VGND VPWR VPWR _1238_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1169_ _2013_/A _2012_/B VGND VGND VPWR VPWR _1170_/B sky130_fd_sc_hd__or2b_2
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2471__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1581__A1 _2409_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2210_ _2204_/Y _2207_/Y _2209_/X VGND VGND VPWR VPWR _2210_/Y sky130_fd_sc_hd__o21ai_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2141_ _2527_/Q VGND VGND VPWR VPWR _2141_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2494__CLK _2512_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2072_ _2294_/A VGND VGND VPWR VPWR _2134_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clkbuf_1_1_0_wb_clk_i/X VGND VGND VPWR VPWR _2576_/CLK sky130_fd_sc_hd__clkbuf_16
X_1925_ _1925_/A VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1856_ _1856_/A VGND VGND VPWR VPWR _1856_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1787_ _2591_/Q _2588_/Q VGND VGND VPWR VPWR _1787_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2408_ _2549_/CLK _2408_/D _1883_/Y VGND VGND VPWR VPWR _2408_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2339_ _2342_/A VGND VGND VPWR VPWR _2339_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1512__B _2028_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input32_A wbs_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ _2397_/Q _2394_/Q VGND VGND VPWR VPWR _1710_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1641_ _2377_/Q _2374_/Q VGND VGND VPWR VPWR _1643_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1572_ input62/X _2413_/Q _1578_/S VGND VGND VPWR VPWR _1573_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2124_ _2117_/Y _2121_/Y _2123_/X VGND VGND VPWR VPWR _2124_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2055_ _1352_/Y _2292_/B _2030_/X _2054_/Y VGND VGND VPWR VPWR _2055_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_78_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1908_ _1912_/A VGND VGND VPWR VPWR _1908_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1839_ _2367_/A VGND VGND VPWR VPWR _1844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2073__B _2134_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput73 _2526_/Q VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput84 _2536_/Q VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput95 _2517_/Q VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2248__B _2285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2255__A2 _2246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2532__CLK _2569_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2264__A _2264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1624_ _2424_/Q VGND VGND VPWR VPWR _1628_/C sky130_fd_sc_hd__inv_2
XFILLER_12_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1555_ _1555_/A VGND VGND VPWR VPWR _2421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1486_ _1486_/A VGND VGND VPWR VPWR _1495_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2107_ _2194_/A _2134_/B _2417_/Q VGND VGND VPWR VPWR _2107_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2038_ _2083_/A _2061_/B _2409_/Q VGND VGND VPWR VPWR _2038_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1489__S _1495_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2182__A1 _2178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2405__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2349__A _2355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2555__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2084__A _2099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ input62/X _1325_/X _1330_/X VGND VGND VPWR VPWR _1340_/X sky130_fd_sc_hd__o21ba_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1271_ _2566_/Q _1261_/X _1267_/X _1270_/Y VGND VGND VPWR VPWR _2565_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2428__CLK _2576_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1607_ _2443_/Q _1586_/B _1596_/X _2445_/Q VGND VGND VPWR VPWR _1608_/C sky130_fd_sc_hd__a31o_1
XFILLER_47_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2587_ _2599_/CLK _2587_/D _2351_/Y VGND VGND VPWR VPWR _2587_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1538_ _1538_/A VGND VGND VPWR VPWR _2429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2578__CLK _2595_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1469_ _2468_/Q _2469_/Q _1473_/S VGND VGND VPWR VPWR _1470_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2510_ _2512_/CLK _2510_/D _2009_/Y VGND VGND VPWR VPWR _2510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2441_ _2599_/CLK _2441_/D _1924_/Y VGND VGND VPWR VPWR _2441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2372_ _2601_/CLK _2372_/D _1838_/Y VGND VGND VPWR VPWR _2372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1323_ _2556_/Q _1311_/X _1317_/X _1322_/Y VGND VGND VPWR VPWR _2555_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1254_ _2568_/Q VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1185_ input6/X input5/X VGND VGND VPWR VPWR _1187_/C sky130_fd_sc_hd__nor2_2
XANTENNA__1621__A _1643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2171__B _2228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input62_A wbs_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1441__A _2448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1941_ _1943_/A VGND VGND VPWR VPWR _1941_/Y sky130_fd_sc_hd__inv_2
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2272__A _2272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1872_ _1875_/A VGND VGND VPWR VPWR _1872_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2424_ _2576_/CLK _2424_/D _1903_/Y VGND VGND VPWR VPWR _2424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2355_ _2355_/A VGND VGND VPWR VPWR _2360_/A sky130_fd_sc_hd__buf_2
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1306_ _2559_/Q _1286_/X _1303_/X _1305_/Y VGND VGND VPWR VPWR _2558_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2286_ _2294_/A _2479_/Q VGND VGND VPWR VPWR _2286_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1237_ _2024_/B VGND VGND VPWR VPWR _1237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1168_ _1165_/Y _1168_/B _1168_/C VGND VGND VPWR VPWR _2014_/A sky130_fd_sc_hd__nand3b_4
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1261__A _1608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2092__A _2099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2133_/Y _2116_/X _2139_/Y VGND VGND VPWR VPWR _2526_/D sky130_fd_sc_hd__o21ai_1
XFILLER_79_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2071_ _2116_/A VGND VGND VPWR VPWR _2071_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1924_ _1925_/A VGND VGND VPWR VPWR _1924_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1855_ _1856_/A VGND VGND VPWR VPWR _1855_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1786_ _2591_/Q _2588_/Q VGND VGND VPWR VPWR _1786_/X sky130_fd_sc_hd__and2_1
XFILLER_102_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2407_ _2459_/CLK _2407_/D _1881_/Y VGND VGND VPWR VPWR _2407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2338_ _2342_/A VGND VGND VPWR VPWR _2338_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2269_ _2263_/Y _2246_/X _2268_/Y VGND VGND VPWR VPWR _2541_/D sky130_fd_sc_hd__o21ai_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2276__B1 _2275_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input25_A wbs_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1640_ _2377_/Q _2374_/Q VGND VGND VPWR VPWR _1643_/D sky130_fd_sc_hd__and2_1
XFILLER_177_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output93_A _2544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1571_ _1571_/A VGND VGND VPWR VPWR _2414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2461__CLK _2549_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_7491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2123_ _2491_/Q _2111_/X _2122_/X _2101_/X VGND VGND VPWR VPWR _2123_/X sky130_fd_sc_hd__o31a_1
XFILLER_3_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2054_ _2054_/A _2452_/Q VGND VGND VPWR VPWR _2054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1907_ _1913_/A VGND VGND VPWR VPWR _1912_/A sky130_fd_sc_hd__buf_2
XFILLER_30_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1838_ _1838_/A VGND VGND VPWR VPWR _1838_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1769_ _1747_/X _2435_/Q _1767_/X _1768_/Y VGND VGND VPWR VPWR _1771_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2484__CLK _2560_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput74 _2527_/Q VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput85 _2537_/Q VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_27_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput96 _2518_/Q VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2264__B _2285_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2278__C_N _2437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1608__B _1608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1623_ _2371_/Q _2368_/Q _1622_/B VGND VGND VPWR VPWR _2371_/D sky130_fd_sc_hd__a21o_1
XFILLER_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1554_ input39/X _2421_/Q _1556_/S VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1485_ _1485_/A VGND VGND VPWR VPWR _2461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

